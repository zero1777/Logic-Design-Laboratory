`define hc  32'd524   // C4
`define hd  32'd588   // D4
`define he  32'd660   // E4
`define hf  32'd698   // F4
`define hg  32'd784   // G4
`define ha  32'd880   // G4
`define hb  32'd988   // G4
`define hhc  32'd1046   // G4
`define da  32'd220   // G4
`define db  32'd245   // G4
`define c   32'd262   // C3
`define d   32'd294   // D3
`define e   32'd330   // D3
`define f   32'd349   // D3
`define g   32'd392   // G3
`define a   32'd440   // G3
`define b   32'd494   // B3
`define rc   32'd277   // c#
`define ld   32'd277   // c#
`define rd   32'd311   // c#
`define le   32'd311   // c#
`define rf   32'd370   // c#
`define lg   32'd370   // c#
`define rg   32'd415   // c#
`define la   32'd415   // c#
`define ra   32'd466   // c#
`define lb   32'd466   // c#
`define rhc   32'd554   // c#
`define lhd   32'd554   // c#
`define rhd   32'd622   // c#
`define lhe   32'd622   // c#
`define rhf   32'd740   // c#
`define lhg   32'd740   // c#
`define rhg   32'd831   // c#
`define lha   32'd831   // c#
`define rha   32'd932   // c#

`define sil   32'd50000000 // slience
`define AA 4'd1
`define BB 4'd2
`define CC 4'd3
`define DD 4'd4
`define EE 4'd5
`define FF 4'd6
`define GG 4'd7


module music_example (
	input [14:0] ibeatNum,
	input en,
    input _music,
	output reg [31:0] toneL,
    output reg [31:0] toneR
);

    always @* begin
        if(en == 1) begin
            if (_music) begin
                case(ibeatNum)
                    // // --- Measure 1 ---
                    // 12'd0: toneR = `hg;      12'd1: toneR = `hg; // HG (half-beat)
                    // 12'd2: toneR = `hg;      12'd3: toneR = `hg;
                    // 12'd4: toneR = `hg;      12'd5: toneR = `hg;
                    // 12'd6: toneR = `hg;      12'd7: toneR = `hg;
                    // 12'd8: toneR = `he;      12'd9: toneR = `he; // HE (half-beat)
                    // 12'd10: toneR = `he;     12'd11: toneR = `he;
                    // 12'd12: toneR = `he;     12'd13: toneR = `he;
                    // 12'd14: toneR = `he;     12'd15: toneR = `sil; // (Short break for repetitive notes: high E)

                    // 12'd16: toneR = `he;     12'd17: toneR = `he; // HE (one-beat)
                    // 12'd18: toneR = `he;     12'd19: toneR = `he;
                    // 12'd20: toneR = `he;     12'd21: toneR = `he;
                    // 12'd22: toneR = `he;     12'd23: toneR = `he;
                    // 12'd24: toneR = `he;     12'd25: toneR = `he;
                    // 12'd26: toneR = `he;     12'd27: toneR = `he;
                    // 12'd28: toneR = `he;     12'd29: toneR = `he;
                    // 12'd30: toneR = `he;     12'd31: toneR = `he;

                    // 12'd32: toneR = `hf;     12'd33: toneR = `hf; // HF (half-beat)
                    // 12'd34: toneR = `hf;     12'd35: toneR = `hf;
                    // 12'd36: toneR = `hf;     12'd37: toneR = `hf;
                    // 12'd38: toneR = `hf;     12'd39: toneR = `hf;
                    // 12'd40: toneR = `hd;     12'd41: toneR = `hd; // HD (half-beat)
                    // 12'd42: toneR = `hd;     12'd43: toneR = `hd;
                    // 12'd44: toneR = `hd;     12'd45: toneR = `hd;
                    // 12'd46: toneR = `hd;     12'd47: toneR = `sil; // (Short break for repetitive notes: high D)

                    // 12'd48: toneR = `hd;     12'd49: toneR = `hd; // HD (one-beat)
                    // 12'd50: toneR = `hd;     12'd51: toneR = `hd;
                    // 12'd52: toneR = `hd;     12'd53: toneR = `hd;
                    // 12'd54: toneR = `hd;     12'd55: toneR = `hd;
                    // 12'd56: toneR = `hd;     12'd57: toneR = `hd;
                    // 12'd58: toneR = `hd;     12'd59: toneR = `hd;
                    // 12'd60: toneR = `hd;     12'd61: toneR = `hd;
                    // 12'd62: toneR = `hd;     12'd63: toneR = `hd;

                    // // --- Measure 2 ---
                    // 12'd64: toneR = `hc;     12'd65: toneR = `hc; // HC (half-beat)
                    // 12'd66: toneR = `hc;     12'd67: toneR = `hc;
                    // 12'd68: toneR = `hc;     12'd69: toneR = `hc;
                    // 12'd70: toneR = `hc;     12'd71: toneR = `hc;
                    // 12'd72: toneR = `hd;     12'd73: toneR = `hd; // HD (half-beat)
                    // 12'd74: toneR = `hd;     12'd75: toneR = `hd;
                    // 12'd76: toneR = `hd;     12'd77: toneR = `hd;
                    // 12'd78: toneR = `hd;     12'd79: toneR = `hd;

                    // 12'd80: toneR = `he;     12'd81: toneR = `he; // HE (half-beat)
                    // 12'd82: toneR = `he;     12'd83: toneR = `he;
                    // 12'd84: toneR = `he;     12'd85: toneR = `he;
                    // 12'd86: toneR = `he;     12'd87: toneR = `he;
                    // 12'd88: toneR = `hf;     12'd89: toneR = `hf; // HF (half-beat)
                    // 12'd90: toneR = `hf;     12'd91: toneR = `hf;
                    // 12'd92: toneR = `hf;     12'd93: toneR = `hf;
                    // 12'd94: toneR = `hf;     12'd95: toneR = `hf;

                    // 12'd96: toneR = `hg;     12'd97: toneR = `hg; // HG (half-beat)
                    // 12'd98: toneR = `hg;     12'd99: toneR = `hg;
                    // 12'd100: toneR = `hg;     12'd101: toneR = `hg;
                    // 12'd102: toneR = `hg;     12'd103: toneR = `sil; // (Short break for repetitive notes: high D)
                    // 12'd104: toneR = `hg;     12'd105: toneR = `hg; // HG (half-beat)
                    // 12'd106: toneR = `hg;     12'd107: toneR = `hg;
                    // 12'd108: toneR = `hg;     12'd109: toneR = `hg;
                    // 12'd110: toneR = `hg;     12'd111: toneR = `sil; // (Short break for repetitive notes: high D)

                    // 12'd112: toneR = `hg;     12'd113: toneR = `hg; // HG (one-beat)
                    // 12'd114: toneR = `hg;     12'd115: toneR = `hg;
                    // 12'd116: toneR = `hg;     12'd117: toneR = `hg;
                    // 12'd118: toneR = `hg;     12'd119: toneR = `hg;
                    // 12'd120: toneR = `hg;     12'd121: toneR = `hg;
                    // 12'd122: toneR = `hg;     12'd123: toneR = `hg;
                    // 12'd124: toneR = `hg;     12'd125: toneR = `hg;
                    // 12'd126: toneR = `hg;     12'd127: toneR = `hg;

                    // 15'd0: toneR = `ha;     15'd1: toneR = `ha;
                    // 15'd2: toneR = `ha;     15'd3: toneR = `ha;
                    // 15'd4: toneR = `ha;     15'd5: toneR = `ha;
                    // 15'd6: toneR = `ha;     15'd7: toneR = `ha;
                    // 15'd8: toneR = `rhf;     15'd9: toneR = `rhf;
                    // 15'd10: toneR = `rhf;     15'd11: toneR = `rhf;
                    // 15'd12: toneR = `hg;     15'd13: toneR = `hg;
                    // 15'd14: toneR = `hg;     15'd15: toneR = `hg;
                    // 15'd16: toneR = `ha;     15'd17: toneR = `ha;
                    // 15'd18: toneR = `ha;     15'd19: toneR = `ha;
                    // 15'd20: toneR = `ha;     15'd21: toneR = `ha;
                    // 15'd22: toneR = `ha;     15'd23: toneR = `ha;
                    // 15'd24: toneR = `rhf;     15'd25: toneR = `rhf;
                    // 15'd26: toneR = `rhf;     15'd27: toneR = `rhf;
                    // 15'd28: toneR = `hg;     15'd29: toneR = `hg;
                    // 15'd30: toneR = `hg;     15'd31: toneR = `hg;
                    // 15'd32: toneR = `ha;     15'd33: toneR = `ha;
                    // 15'd34: toneR = `ha;     15'd35: toneR = `ha;
                    // 15'd36: toneR = `a;     15'd37: toneR = `a;
                    // 15'd38: toneR = `a;     15'd39: toneR = `a;
                    // 15'd40: toneR = `b;     15'd41: toneR = `b;
                    // 15'd42: toneR = `b;     15'd43: toneR = `b;
                    // 15'd44: toneR = `rhc;     15'd45: toneR = `rhc;
                    // 15'd46: toneR = `rhc;     15'd47: toneR = `rhc;
                    // 15'd48: toneR = `hd;     15'd49: toneR = `hd;
                    // 15'd50: toneR = `hd;     15'd51: toneR = `hd;
                    // 15'd52: toneR = `he;     15'd53: toneR = `he;
                    // 15'd54: toneR = `he;     15'd55: toneR = `he;
                    // 15'd56: toneR = `rhf;     15'd57: toneR = `rhf;
                    // 15'd58: toneR = `rhf;     15'd59: toneR = `rhf;
                    // 15'd60: toneR = `hg;     15'd61: toneR = `hg;
                    // 15'd62: toneR = `hg;     15'd63: toneR = `hg;
                    // 15'd64: toneR = `rhf;     15'd65: toneR = `rhf;
                    // 15'd66: toneR = `rhf;     15'd67: toneR = `rhf;
                    // 15'd68: toneR = `rhf;     15'd69: toneR = `rhf;
                    // 15'd70: toneR = `rhf;     15'd71: toneR = `rhf;
                    // 15'd72: toneR = `hd;     15'd73: toneR = `hd;
                    // 15'd74: toneR = `hd;     15'd75: toneR = `hd;
                    // 15'd76: toneR = `he;     15'd77: toneR = `he;
                    // 15'd78: toneR = `he;     15'd79: toneR = `he;
                    // 15'd80: toneR = `rhf;     15'd81: toneR = `rhf;
                    // 15'd82: toneR = `rhf;     15'd83: toneR = `rhf;
                    // 15'd84: toneR = `rhf;     15'd85: toneR = `rhf;
                    // 15'd86: toneR = `rhf;     15'd87: toneR = `rhf;
                    // 15'd88: toneR = `rf;     15'd89: toneR = `rf;
                    // 15'd90: toneR = `rf;     15'd91: toneR = `rf;
                    // 15'd92: toneR = `g;     15'd93: toneR = `g;
                    // 15'd94: toneR = `g;     15'd95: toneR = `g;
                    // 15'd96: toneR = `a;     15'd97: toneR = `a;
                    // 15'd98: toneR = `a;     15'd99: toneR = `a;
                    // 15'd100: toneR = `b;     15'd101: toneR = `b;
                    // 15'd102: toneR = `b;     15'd103: toneR = `b;
                    // 15'd104: toneR = `a;     15'd105: toneR = `a;
                    // 15'd106: toneR = `a;     15'd107: toneR = `a;
                    // 15'd108: toneR = `g;     15'd109: toneR = `g;
                    // 15'd110: toneR = `g;     15'd111: toneR = `g;
                    // 15'd112: toneR = `a;     15'd113: toneR = `a;
                    // 15'd114: toneR = `a;     15'd115: toneR = `a;
                    // 15'd116: toneR = `rf;     15'd117: toneR = `rf;
                    // 15'd118: toneR = `rf;     15'd119: toneR = `rf;
                    // 15'd120: toneR = `g;     15'd121: toneR = `g;
                    // 15'd122: toneR = `g;     15'd123: toneR = `g;
                    // 15'd124: toneR = `a;     15'd125: toneR = `a;
                    // 15'd126: toneR = `a;     15'd127: toneR = `a;
                    // 15'd128: toneR = `g;     15'd129: toneR = `g;
                    // 15'd130: toneR = `g;     15'd131: toneR = `g;
                    // 15'd132: toneR = `g;     15'd133: toneR = `g;
                    // 15'd134: toneR = `g;     15'd135: toneR = `g;
                    // 15'd136: toneR = `b;     15'd137: toneR = `b;
                    // 15'd138: toneR = `b;     15'd139: toneR = `b;
                    // 15'd140: toneR = `a;     15'd141: toneR = `a;
                    // 15'd142: toneR = `a;     15'd143: toneR = `a;
                    // 15'd144: toneR = `g;     15'd145: toneR = `g;
                    // 15'd146: toneR = `g;     15'd147: toneR = `g;
                    // 15'd148: toneR = `g;     15'd149: toneR = `g;
                    // 15'd150: toneR = `g;     15'd151: toneR = `g;
                    // 15'd152: toneR = `rf;     15'd153: toneR = `rf;
                    // 15'd154: toneR = `rf;     15'd155: toneR = `rf;
                    // 15'd156: toneR = `e;     15'd157: toneR = `e;
                    // 15'd158: toneR = `e;     15'd159: toneR = `e;
                    // 15'd160: toneR = `rf;     15'd161: toneR = `rf;
                    // 15'd162: toneR = `rf;     15'd163: toneR = `rf;
                    // 15'd164: toneR = `e;     15'd165: toneR = `e;
                    // 15'd166: toneR = `e;     15'd167: toneR = `e;
                    // 15'd168: toneR = `d;     15'd169: toneR = `d;
                    // 15'd170: toneR = `d;     15'd171: toneR = `d;
                    // 15'd172: toneR = `e;     15'd173: toneR = `e;
                    // 15'd174: toneR = `e;     15'd175: toneR = `e;
                    // 15'd176: toneR = `rf;     15'd177: toneR = `rf;
                    // 15'd178: toneR = `rf;     15'd179: toneR = `rf;
                    // 15'd180: toneR = `g;     15'd181: toneR = `g;
                    // 15'd182: toneR = `g;     15'd183: toneR = `g;
                    // 15'd184: toneR = `a;     15'd185: toneR = `a;
                    // 15'd186: toneR = `a;     15'd187: toneR = `a;
                    // 15'd188: toneR = `b;     15'd189: toneR = `b;
                    // 15'd190: toneR = `b;     15'd191: toneR = `b;
                    // 15'd192: toneR = `g;     15'd193: toneR = `g;
                    // 15'd194: toneR = `g;     15'd195: toneR = `g;
                    // 15'd196: toneR = `g;     15'd197: toneR = `g;
                    // 15'd198: toneR = `g;     15'd199: toneR = `g;
                    // 15'd200: toneR = `b;     15'd201: toneR = `b;
                    // 15'd202: toneR = `b;     15'd203: toneR = `b;
                    // 15'd204: toneR = `a;     15'd205: toneR = `a;
                    // 15'd206: toneR = `a;     15'd207: toneR = `a;
                    // 15'd208: toneR = `b;     15'd209: toneR = `b;
                    // 15'd210: toneR = `b;     15'd211: toneR = `b;
                    // 15'd212: toneR = `b;     15'd213: toneR = `b;
                    // 15'd214: toneR = `b;     15'd215: toneR = `b;
                    // 15'd216: toneR = `rhc;     15'd217: toneR = `rhc;
                    // 15'd218: toneR = `rhc;     15'd219: toneR = `rhc;
                    // 15'd220: toneR = `hd;     15'd221: toneR = `hd;
                    // 15'd222: toneR = `hd;     15'd223: toneR = `hd;
                    // 15'd224: toneR = `a;     15'd225: toneR = `a;
                    // 15'd226: toneR = `a;     15'd227: toneR = `a;
                    // 15'd228: toneR = `b;     15'd229: toneR = `b;
                    // 15'd230: toneR = `b;     15'd231: toneR = `b;
                    // 15'd232: toneR = `rhc;     15'd233: toneR = `rhc;
                    // 15'd234: toneR = `rhc;     15'd235: toneR = `rhc;
                    // 15'd236: toneR = `hd;     15'd237: toneR = `hd;
                    // 15'd238: toneR = `hd;     15'd239: toneR = `hd;
                    // 15'd240: toneR = `he;     15'd241: toneR = `he;
                    // 15'd242: toneR = `he;     15'd243: toneR = `he;
                    // 15'd244: toneR = `rhf;     15'd245: toneR = `rhf;
                    // 15'd246: toneR = `rhf;     15'd247: toneR = `rhf;
                    // 15'd248: toneR = `hg;     15'd249: toneR = `hg;
                    // 15'd250: toneR = `hg;     15'd251: toneR = `hg;
                    // 15'd252: toneR = `ha;     15'd253: toneR = `ha;
                    // 15'd254: toneR = `ha;     15'd255: toneR = `ha;
                    // 15'd256: toneR = `rhf;     15'd257: toneR = `rhf;
                    // 15'd258: toneR = `rhf;     15'd259: toneR = `rhf;
                    // 15'd260: toneR = `rhf;     15'd261: toneR = `rhf;
                    // 15'd262: toneR = `rhf;     15'd263: toneR = `rhf;
                    // 15'd264: toneR = `hd;     15'd265: toneR = `hd;
                    // 15'd266: toneR = `hd;     15'd267: toneR = `hd;
                    // 15'd268: toneR = `he;     15'd269: toneR = `he;
                    // 15'd270: toneR = `he;     15'd271: toneR = `he;
                    // 15'd272: toneR = `rhf;     15'd273: toneR = `rhf;
                    // 15'd274: toneR = `rhf;     15'd275: toneR = `rhf;
                    // 15'd276: toneR = `rhf;     15'd277: toneR = `rhf;
                    // 15'd278: toneR = `rhf;     15'd279: toneR = `rhf;
                    // 15'd280: toneR = `he;     15'd281: toneR = `he;
                    // 15'd282: toneR = `he;     15'd283: toneR = `he;
                    // 15'd284: toneR = `hd;     15'd285: toneR = `hd;
                    // 15'd286: toneR = `hd;     15'd287: toneR = `hd;
                    // 15'd288: toneR = `he;     15'd289: toneR = `he;
                    // 15'd290: toneR = `he;     15'd291: toneR = `he;
                    // 15'd292: toneR = `rhc;     15'd293: toneR = `rhc;
                    // 15'd294: toneR = `rhc;     15'd295: toneR = `rhc;
                    // 15'd296: toneR = `hd;     15'd297: toneR = `hd;
                    // 15'd298: toneR = `hd;     15'd299: toneR = `hd;
                    // 15'd300: toneR = `he;     15'd301: toneR = `he;
                    // 15'd302: toneR = `he;     15'd303: toneR = `he;
                    // 15'd304: toneR = `rhf;     15'd305: toneR = `rhf;
                    // 15'd306: toneR = `rhf;     15'd307: toneR = `rhf;
                    // 15'd308: toneR = `he;     15'd309: toneR = `he;
                    // 15'd310: toneR = `he;     15'd311: toneR = `he;
                    // 15'd312: toneR = `hd;     15'd313: toneR = `hd;
                    // 15'd314: toneR = `hd;     15'd315: toneR = `hd;
                    // 15'd316: toneR = `rhc;     15'd317: toneR = `rhc;
                    // 15'd318: toneR = `rhc;     15'd319: toneR = `rhc;

                    15'd0: toneR = `e;     15'd1: toneR = `e;
15'd2: toneR = `e;     15'd3: toneR = `e;
15'd4: toneR = `f;     15'd5: toneR = `f;
15'd6: toneR = `f;     15'd7: toneR = `f;
15'd8: toneR = `g;     15'd9: toneR = `g;
15'd10: toneR = `g;     15'd11: toneR = `g;
15'd12: toneR = `g;     15'd13: toneR = `g;
15'd14: toneR = `g;     15'd15: toneR = `g;
15'd16: toneR = `g;     15'd17: toneR = `g;
15'd18: toneR = `g;     15'd19: toneR = `g;
15'd20: toneR = `g;     15'd21: toneR = `g;
15'd22: toneR = `g;     15'd23: toneR = `g;
15'd24: toneR = `sil;     15'd25: toneR = `g;
15'd26: toneR = `g;     15'd27: toneR = `g;
15'd28: toneR = `g;     15'd29: toneR = `g;
15'd30: toneR = `g;     15'd31: toneR = `g;
15'd32: toneR = `g;     15'd33: toneR = `g;
15'd34: toneR = `g;     15'd35: toneR = `g;
15'd36: toneR = `g;     15'd37: toneR = `g;
15'd38: toneR = `g;     15'd39: toneR = `g;
15'd40: toneR = `f;     15'd41: toneR = `f;
15'd42: toneR = `f;     15'd43: toneR = `f;
15'd44: toneR = `f;     15'd45: toneR = `f;
15'd46: toneR = `f;     15'd47: toneR = `f;
15'd48: toneR = `e;     15'd49: toneR = `e;
15'd50: toneR = `e;     15'd51: toneR = `e;
15'd52: toneR = `e;     15'd53: toneR = `e;
15'd54: toneR = `e;     15'd55: toneR = `e;
15'd56: toneR = `d;     15'd57: toneR = `d;
15'd58: toneR = `d;     15'd59: toneR = `d;
15'd60: toneR = `d;     15'd61: toneR = `d;
15'd62: toneR = `d;     15'd63: toneR = `d;
15'd64: toneR = `c;     15'd65: toneR = `c;
15'd66: toneR = `c;     15'd67: toneR = `c;
15'd68: toneR = `c;     15'd69: toneR = `c;
15'd70: toneR = `c;     15'd71: toneR = `c;
15'd72: toneR = `db;     15'd73: toneR = `db;
15'd74: toneR = `db;     15'd75: toneR = `db;
15'd76: toneR = `db;     15'd77: toneR = `db;
15'd78: toneR = `db;     15'd79: toneR = `db;
15'd80: toneR = `g;     15'd81: toneR = `g;
15'd82: toneR = `g;     15'd83: toneR = `g;
15'd84: toneR = `g;     15'd85: toneR = `g;
15'd86: toneR = `g;     15'd87: toneR = `g;
15'd88: toneR = `g;     15'd89: toneR = `g;
15'd90: toneR = `g;     15'd91: toneR = `g;
15'd92: toneR = `g;     15'd93: toneR = `g;
15'd94: toneR = `g;     15'd95: toneR = `g;
15'd96: toneR = `e;     15'd97: toneR = `e;
15'd98: toneR = `e;     15'd99: toneR = `e;
15'd100: toneR = `e;     15'd101: toneR = `e;
15'd102: toneR = `e;     15'd103: toneR = `e;
15'd104: toneR = `e;     15'd105: toneR = `e;
15'd106: toneR = `e;     15'd107: toneR = `e;
15'd108: toneR = `e;     15'd109: toneR = `e;
15'd110: toneR = `e;     15'd111: toneR = `e;
15'd112: toneR = `e;     15'd113: toneR = `e;
15'd114: toneR = `e;     15'd115: toneR = `e;
15'd116: toneR = `e;     15'd117: toneR = `e;
15'd118: toneR = `e;     15'd119: toneR = `e;
15'd120: toneR = `e;     15'd121: toneR = `e;
15'd122: toneR = `e;     15'd123: toneR = `e;
15'd124: toneR = `e;     15'd125: toneR = `e;
15'd126: toneR = `e;     15'd127: toneR = `e;
15'd128: toneR = `e;     15'd129: toneR = `e;
15'd130: toneR = `e;     15'd131: toneR = `e;
15'd132: toneR = `e;     15'd133: toneR = `e;
15'd134: toneR = `e;     15'd135: toneR = `e;
15'd136: toneR = `c;     15'd137: toneR = `c;
15'd138: toneR = `c;     15'd139: toneR = `c;
15'd140: toneR = `c;     15'd141: toneR = `c;
15'd142: toneR = `c;     15'd143: toneR = `c;
15'd144: toneR = `c;     15'd145: toneR = `c;
15'd146: toneR = `c;     15'd147: toneR = `c;
15'd148: toneR = `c;     15'd149: toneR = `c;
15'd150: toneR = `c;     15'd151: toneR = `c;
15'd152: toneR = `g;     15'd153: toneR = `g;
15'd154: toneR = `g;     15'd155: toneR = `g;
15'd156: toneR = `g;     15'd157: toneR = `g;
15'd158: toneR = `g;     15'd159: toneR = `g;
15'd160: toneR = `g;     15'd161: toneR = `g;
15'd162: toneR = `g;     15'd163: toneR = `g;
15'd164: toneR = `g;     15'd165: toneR = `g;
15'd166: toneR = `g;     15'd167: toneR = `g;
15'd168: toneR = `f;     15'd169: toneR = `f;
15'd170: toneR = `f;     15'd171: toneR = `f;
15'd172: toneR = `f;     15'd173: toneR = `f;
15'd174: toneR = `f;     15'd175: toneR = `f;
15'd176: toneR = `e;     15'd177: toneR = `e;
15'd178: toneR = `e;     15'd179: toneR = `e;
15'd180: toneR = `e;     15'd181: toneR = `e;
15'd182: toneR = `e;     15'd183: toneR = `e;
15'd184: toneR = `d;     15'd185: toneR = `d;
15'd186: toneR = `d;     15'd187: toneR = `d;
15'd188: toneR = `d;     15'd189: toneR = `d;
15'd190: toneR = `d;     15'd191: toneR = `d;
15'd192: toneR = `c;     15'd193: toneR = `c;
15'd194: toneR = `c;     15'd195: toneR = `c;
15'd196: toneR = `c;     15'd197: toneR = `c;
15'd198: toneR = `c;     15'd199: toneR = `c;
15'd200: toneR = `d;     15'd201: toneR = `d;
15'd202: toneR = `d;     15'd203: toneR = `d;
15'd204: toneR = `d;     15'd205: toneR = `d;
15'd206: toneR = `d;     15'd207: toneR = `d;
15'd208: toneR = `d;     15'd209: toneR = `d;
15'd210: toneR = `d;     15'd211: toneR = `d;
15'd212: toneR = `d;     15'd213: toneR = `d;
15'd214: toneR = `d;     15'd215: toneR = `d;
15'd216: toneR = `d;     15'd217: toneR = `d;
15'd218: toneR = `d;     15'd219: toneR = `d;
15'd220: toneR = `d;     15'd221: toneR = `d;
15'd222: toneR = `d;     15'd223: toneR = `d;
15'd224: toneR = `c;     15'd225: toneR = `c;
15'd226: toneR = `c;     15'd227: toneR = `c;
15'd228: toneR = `c;     15'd229: toneR = `c;
15'd230: toneR = `c;     15'd231: toneR = `c;
15'd232: toneR = `sil;     15'd233: toneR = `c;
15'd234: toneR = `c;     15'd235: toneR = `c;
15'd236: toneR = `c;     15'd237: toneR = `c;
15'd238: toneR = `c;     15'd239: toneR = `c;
15'd240: toneR = `c;     15'd241: toneR = `c;
15'd242: toneR = `c;     15'd243: toneR = `c;
15'd244: toneR = `c;     15'd245: toneR = `c;
15'd246: toneR = `c;     15'd247: toneR = `c;
15'd248: toneR = `sil;     15'd249: toneR = `sil;
15'd250: toneR = `sil;     15'd251: toneR = `sil;
15'd252: toneR = `sil;     15'd253: toneR = `sil;
15'd254: toneR = `sil;     15'd255: toneR = `sil;
15'd256: toneR = `e;     15'd257: toneR = `e;
15'd258: toneR = `e;     15'd259: toneR = `e;
15'd260: toneR = `f;     15'd261: toneR = `f;
15'd262: toneR = `f;     15'd263: toneR = `f;
15'd264: toneR = `g;     15'd265: toneR = `g;
15'd266: toneR = `g;     15'd267: toneR = `g;
15'd268: toneR = `g;     15'd269: toneR = `g;
15'd270: toneR = `g;     15'd271: toneR = `g;
15'd272: toneR = `sil;     15'd273: toneR = `g;
15'd274: toneR = `g;     15'd275: toneR = `g;
15'd276: toneR = `g;     15'd277: toneR = `g;
15'd278: toneR = `g;     15'd279: toneR = `g;
15'd280: toneR = `sil;     15'd281: toneR = `g;
15'd282: toneR = `g;     15'd283: toneR = `g;
15'd284: toneR = `g;     15'd285: toneR = `g;
15'd286: toneR = `a;     15'd287: toneR = `a;
15'd288: toneR = `a;     15'd289: toneR = `a;
15'd290: toneR = `a;     15'd291: toneR = `a;
15'd292: toneR = `a;     15'd293: toneR = `a;
15'd294: toneR = `a;     15'd295: toneR = `a;
15'd296: toneR = `g;     15'd297: toneR = `g;
15'd298: toneR = `g;     15'd299: toneR = `g;
15'd300: toneR = `g;     15'd301: toneR = `g;
15'd302: toneR = `g;     15'd303: toneR = `g;
15'd304: toneR = `g;     15'd305: toneR = `g;
15'd306: toneR = `g;     15'd307: toneR = `g;
15'd308: toneR = `g;     15'd309: toneR = `g;
15'd310: toneR = `g;     15'd311: toneR = `g;
15'd312: toneR = `g;     15'd313: toneR = `g;
15'd314: toneR = `g;     15'd315: toneR = `g;
15'd316: toneR = `g;     15'd317: toneR = `g;
15'd318: toneR = `g;     15'd319: toneR = `g;
15'd320: toneR = `e;     15'd321: toneR = `e;
15'd322: toneR = `e;     15'd323: toneR = `e;
15'd324: toneR = `f;     15'd325: toneR = `f;
15'd326: toneR = `f;     15'd327: toneR = `f;
15'd328: toneR = `g;     15'd329: toneR = `g;
15'd330: toneR = `g;     15'd331: toneR = `g;
15'd332: toneR = `g;     15'd333: toneR = `g;
15'd334: toneR = `g;     15'd335: toneR = `g;
15'd336: toneR = `sil;     15'd337: toneR = `g;
15'd338: toneR = `g;     15'd339: toneR = `g;
15'd340: toneR = `g;     15'd341: toneR = `g;
15'd342: toneR = `g;     15'd343: toneR = `g;
15'd344: toneR = `sil;     15'd345: toneR = `g;
15'd346: toneR = `g;     15'd347: toneR = `g;
15'd348: toneR = `g;     15'd349: toneR = `g;
15'd350: toneR = `g;     15'd351: toneR = `g;
15'd352: toneR = `d;     15'd353: toneR = `d;
15'd354: toneR = `d;     15'd355: toneR = `d;
15'd356: toneR = `d;     15'd357: toneR = `d;
15'd358: toneR = `d;     15'd359: toneR = `d;
15'd360: toneR = `e;     15'd361: toneR = `e;
15'd362: toneR = `e;     15'd363: toneR = `e;
15'd364: toneR = `e;     15'd365: toneR = `e;
15'd366: toneR = `e;     15'd367: toneR = `e;
15'd368: toneR = `e;     15'd369: toneR = `e;
15'd370: toneR = `e;     15'd371: toneR = `e;
15'd372: toneR = `e;     15'd373: toneR = `e;
15'd374: toneR = `e;     15'd375: toneR = `e;
15'd376: toneR = `e;     15'd377: toneR = `e;
15'd378: toneR = `e;     15'd379: toneR = `e;
15'd380: toneR = `e;     15'd381: toneR = `e;
15'd382: toneR = `e;     15'd383: toneR = `e;
15'd384: toneR = `sil;     15'd385: toneR = `e;
15'd386: toneR = `e;     15'd387: toneR = `e;
15'd388: toneR = `f;     15'd389: toneR = `f;
15'd390: toneR = `f;     15'd391: toneR = `f;
15'd392: toneR = `g;     15'd393: toneR = `g;
15'd394: toneR = `g;     15'd395: toneR = `g;
15'd396: toneR = `g;     15'd397: toneR = `g;
15'd398: toneR = `g;     15'd399: toneR = `g;
15'd400: toneR = `sil;     15'd401: toneR = `g;
15'd402: toneR = `g;     15'd403: toneR = `g;
15'd404: toneR = `sil;     15'd405: toneR = `g;
15'd406: toneR = `g;     15'd407: toneR = `g;
15'd408: toneR = `g;     15'd409: toneR = `g;
15'd410: toneR = `g;     15'd411: toneR = `g;
15'd412: toneR = `g;     15'd413: toneR = `g;
15'd414: toneR = `sil;     15'd415: toneR = `g;
15'd416: toneR = `g;     15'd417: toneR = `g;
15'd418: toneR = `g;     15'd419: toneR = `g;
15'd420: toneR = `g;     15'd421: toneR = `g;
15'd422: toneR = `sil;     15'd423: toneR = `sil;
15'd424: toneR = `a;     15'd425: toneR = `a;
15'd426: toneR = `a;     15'd427: toneR = `a;
15'd428: toneR = `a;     15'd429: toneR = `a;
15'd430: toneR = `a;     15'd431: toneR = `a;
15'd432: toneR = `g;     15'd433: toneR = `g;
15'd434: toneR = `g;     15'd435: toneR = `g;
15'd436: toneR = `g;     15'd437: toneR = `g;
15'd438: toneR = `g;     15'd439: toneR = `g;
15'd440: toneR = `f;     15'd441: toneR = `f;
15'd442: toneR = `f;     15'd443: toneR = `f;
15'd444: toneR = `f;     15'd445: toneR = `f;
15'd446: toneR = `f;     15'd447: toneR = `f;
15'd448: toneR = `e;     15'd449: toneR = `e;
15'd450: toneR = `e;     15'd451: toneR = `e;
15'd452: toneR = `e;     15'd453: toneR = `e;
15'd454: toneR = `e;     15'd455: toneR = `e;
15'd456: toneR = `d;     15'd457: toneR = `d;
15'd458: toneR = `d;     15'd459: toneR = `d;
15'd460: toneR = `d;     15'd461: toneR = `d;
15'd462: toneR = `d;     15'd463: toneR = `d;
15'd464: toneR = `d;     15'd465: toneR = `d;
15'd466: toneR = `d;     15'd467: toneR = `d;
15'd468: toneR = `d;     15'd469: toneR = `d;
15'd470: toneR = `d;     15'd471: toneR = `d;
15'd472: toneR = `e;     15'd473: toneR = `e;
15'd474: toneR = `e;     15'd475: toneR = `e;
15'd476: toneR = `e;     15'd477: toneR = `e;
15'd478: toneR = `e;     15'd479: toneR = `e;
15'd480: toneR = `e;     15'd481: toneR = `e;
15'd482: toneR = `e;     15'd483: toneR = `e;
15'd484: toneR = `e;     15'd485: toneR = `e;
15'd486: toneR = `e;     15'd487: toneR = `e;
15'd488: toneR = `sil;     15'd489: toneR = `e;
15'd490: toneR = `e;     15'd491: toneR = `e;
15'd492: toneR = `e;     15'd493: toneR = `e;
15'd494: toneR = `e;     15'd495: toneR = `e;
15'd496: toneR = `e;     15'd497: toneR = `e;
15'd498: toneR = `e;     15'd499: toneR = `e;
15'd500: toneR = `e;     15'd501: toneR = `e;
15'd502: toneR = `e;     15'd503: toneR = `e;
15'd504: toneR = `hc;     15'd505: toneR = `hc;
15'd506: toneR = `hc;     15'd507: toneR = `hc;
15'd508: toneR = `hc;     15'd509: toneR = `hc;
15'd510: toneR = `hc;     15'd511: toneR = `hc;
15'd512: toneR = `b;     15'd513: toneR = `b;
15'd514: toneR = `b;     15'd515: toneR = `b;
15'd516: toneR = `b;     15'd517: toneR = `b;
15'd518: toneR = `b;     15'd519: toneR = `b;
15'd520: toneR = `a;     15'd521: toneR = `a;
15'd522: toneR = `a;     15'd523: toneR = `a;
15'd524: toneR = `a;     15'd525: toneR = `a;
15'd526: toneR = `a;     15'd527: toneR = `a;
15'd528: toneR = `g;     15'd529: toneR = `g;
15'd530: toneR = `g;     15'd531: toneR = `g;
15'd532: toneR = `g;     15'd533: toneR = `g;
15'd534: toneR = `g;     15'd535: toneR = `g;
15'd536: toneR = `e;     15'd537: toneR = `e;
15'd538: toneR = `e;     15'd539: toneR = `e;
15'd540: toneR = `e;     15'd541: toneR = `e;
15'd542: toneR = `e;     15'd543: toneR = `e;
15'd544: toneR = `d;     15'd545: toneR = `d;
15'd546: toneR = `d;     15'd547: toneR = `d;
15'd548: toneR = `sil;     15'd549: toneR = `d;
15'd550: toneR = `d;     15'd551: toneR = `d;
15'd552: toneR = `d;     15'd553: toneR = `d;
15'd554: toneR = `d;     15'd555: toneR = `d;
15'd556: toneR = `d;     15'd557: toneR = `d;
15'd558: toneR = `d;     15'd559: toneR = `d;
15'd560: toneR = `c;     15'd561: toneR = `c;
15'd562: toneR = `c;     15'd563: toneR = `c;
15'd564: toneR = `c;     15'd565: toneR = `c;
15'd566: toneR = `c;     15'd567: toneR = `c;
15'd568: toneR = `da;     15'd569: toneR = `da;
15'd570: toneR = `da;     15'd571: toneR = `da;
15'd572: toneR = `da;     15'd573: toneR = `da;
15'd574: toneR = `da;     15'd575: toneR = `da;
15'd576: toneR = `db;     15'd577: toneR = `db;
15'd578: toneR = `db;     15'd579: toneR = `db;
15'd580: toneR = `c;     15'd581: toneR = `c;
15'd582: toneR = `c;     15'd583: toneR = `c;
15'd584: toneR = `c;     15'd585: toneR = `c;
15'd586: toneR = `c;     15'd587: toneR = `c;
15'd588: toneR = `c;     15'd589: toneR = `c;
15'd590: toneR = `c;     15'd591: toneR = `c;
15'd592: toneR = `c;     15'd593: toneR = `c;
15'd594: toneR = `c;     15'd595: toneR = `c;
15'd596: toneR = `c;     15'd597: toneR = `c;
15'd598: toneR = `c;     15'd599: toneR = `c;
15'd600: toneR = `sil;     15'd601: toneR = `sil;
15'd602: toneR = `sil;     15'd603: toneR = `sil;
15'd604: toneR = `sil;     15'd605: toneR = `sil;
15'd606: toneR = `sil;     15'd607: toneR = `sil;
15'd608: toneR = `sil;     15'd609: toneR = `sil;
15'd610: toneR = `sil;     15'd611: toneR = `sil;
15'd612: toneR = `sil;     15'd613: toneR = `sil;
15'd614: toneR = `sil;     15'd615: toneR = `sil;
15'd616: toneR = `sil;     15'd617: toneR = `sil;
15'd618: toneR = `sil;     15'd619: toneR = `sil;
15'd620: toneR = `sil;     15'd621: toneR = `sil;
15'd622: toneR = `sil;     15'd623: toneR = `sil;
15'd624: toneR = `sil;     15'd625: toneR = `sil;
15'd626: toneR = `sil;     15'd627: toneR = `sil;
15'd628: toneR = `sil;     15'd629: toneR = `sil;
15'd630: toneR = `sil;     15'd631: toneR = `sil;
15'd632: toneR = `sil;     15'd633: toneR = `sil;
15'd634: toneR = `sil;     15'd635: toneR = `sil;
15'd636: toneR = `sil;     15'd637: toneR = `sil;
15'd638: toneR = `sil;     15'd639: toneR = `sil;
15'd640: toneR = `sil;     15'd641: toneR = `sil;
15'd642: toneR = `sil;     15'd643: toneR = `sil;
15'd644: toneR = `sil;     15'd645: toneR = `sil;
15'd646: toneR = `sil;     15'd647: toneR = `sil;
15'd648: toneR = `sil;     15'd649: toneR = `sil;
15'd650: toneR = `sil;     15'd651: toneR = `sil;
15'd652: toneR = `sil;     15'd653: toneR = `sil;
15'd654: toneR = `sil;     15'd655: toneR = `sil;
15'd656: toneR = `sil;     15'd657: toneR = `sil;
15'd658: toneR = `sil;     15'd659: toneR = `sil;
15'd660: toneR = `sil;     15'd661: toneR = `sil;
15'd662: toneR = `sil;     15'd663: toneR = `sil;
15'd664: toneR = `sil;     15'd665: toneR = `sil;
15'd666: toneR = `sil;     15'd667: toneR = `sil;
15'd668: toneR = `sil;     15'd669: toneR = `sil;
15'd670: toneR = `sil;     15'd671: toneR = `sil;
15'd672: toneR = `sil;     15'd673: toneR = `sil;
15'd674: toneR = `sil;     15'd675: toneR = `sil;
15'd676: toneR = `sil;     15'd677: toneR = `sil;
15'd678: toneR = `sil;     15'd679: toneR = `sil;
15'd680: toneR = `sil;     15'd681: toneR = `sil;
15'd682: toneR = `sil;     15'd683: toneR = `sil;
15'd684: toneR = `sil;     15'd685: toneR = `sil;
15'd686: toneR = `sil;     15'd687: toneR = `sil;
15'd688: toneR = `sil;     15'd689: toneR = `sil;
15'd690: toneR = `sil;     15'd691: toneR = `sil;
15'd692: toneR = `sil;     15'd693: toneR = `sil;
15'd694: toneR = `sil;     15'd695: toneR = `sil;
15'd696: toneR = `sil;     15'd697: toneR = `sil;
15'd698: toneR = `sil;     15'd699: toneR = `sil;
15'd700: toneR = `sil;     15'd701: toneR = `sil;
15'd702: toneR = `sil;     15'd703: toneR = `sil;
15'd704: toneR = `e;     15'd705: toneR = `e;
15'd706: toneR = `e;     15'd707: toneR = `e;
15'd708: toneR = `f;     15'd709: toneR = `f;
15'd710: toneR = `f;     15'd711: toneR = `f;
15'd712: toneR = `g;     15'd713: toneR = `g;
15'd714: toneR = `g;     15'd715: toneR = `g;
15'd716: toneR = `g;     15'd717: toneR = `g;
15'd718: toneR = `g;     15'd719: toneR = `g;
15'd720: toneR = `sil;     15'd721: toneR = `g;
15'd722: toneR = `g;     15'd723: toneR = `g;
15'd724: toneR = `g;     15'd725: toneR = `g;
15'd726: toneR = `g;     15'd727: toneR = `g;
15'd728: toneR = `sil;     15'd729: toneR = `g;
15'd730: toneR = `g;     15'd731: toneR = `g;
15'd732: toneR = `g;     15'd733: toneR = `g;
15'd734: toneR = `a;     15'd735: toneR = `a;
15'd736: toneR = `a;     15'd737: toneR = `a;
15'd738: toneR = `a;     15'd739: toneR = `a;
15'd740: toneR = `a;     15'd741: toneR = `a;
15'd742: toneR = `a;     15'd743: toneR = `a;
15'd744: toneR = `g;     15'd745: toneR = `g;
15'd746: toneR = `g;     15'd747: toneR = `g;
15'd748: toneR = `g;     15'd749: toneR = `g;
15'd750: toneR = `g;     15'd751: toneR = `g;
15'd752: toneR = `g;     15'd753: toneR = `g;
15'd754: toneR = `g;     15'd755: toneR = `g;
15'd756: toneR = `g;     15'd757: toneR = `g;
15'd758: toneR = `g;     15'd759: toneR = `g;
15'd760: toneR = `g;     15'd761: toneR = `g;
15'd762: toneR = `g;     15'd763: toneR = `g;
15'd764: toneR = `g;     15'd765: toneR = `g;
15'd766: toneR = `g;     15'd767: toneR = `g;
15'd768: toneR = `e;     15'd769: toneR = `e;
15'd770: toneR = `e;     15'd771: toneR = `e;
15'd772: toneR = `f;     15'd773: toneR = `f;
15'd774: toneR = `f;     15'd775: toneR = `f;
15'd776: toneR = `g;     15'd777: toneR = `g;
15'd778: toneR = `g;     15'd779: toneR = `g;
15'd780: toneR = `g;     15'd781: toneR = `g;
15'd782: toneR = `g;     15'd783: toneR = `g;
15'd784: toneR = `sil;     15'd785: toneR = `g;
15'd786: toneR = `g;     15'd787: toneR = `g;
15'd788: toneR = `g;     15'd789: toneR = `g;
15'd790: toneR = `g;     15'd791: toneR = `g;
15'd792: toneR = `sil;     15'd793: toneR = `g;
15'd794: toneR = `g;     15'd795: toneR = `g;
15'd796: toneR = `g;     15'd797: toneR = `g;
15'd798: toneR = `g;     15'd799: toneR = `g;
15'd800: toneR = `d;     15'd801: toneR = `d;
15'd802: toneR = `d;     15'd803: toneR = `d;
15'd804: toneR = `d;     15'd805: toneR = `d;
15'd806: toneR = `d;     15'd807: toneR = `d;
15'd808: toneR = `e;     15'd809: toneR = `e;
15'd810: toneR = `e;     15'd811: toneR = `e;
15'd812: toneR = `e;     15'd813: toneR = `e;
15'd814: toneR = `e;     15'd815: toneR = `e;
15'd816: toneR = `e;     15'd817: toneR = `e;
15'd818: toneR = `e;     15'd819: toneR = `e;
15'd820: toneR = `e;     15'd821: toneR = `e;
15'd822: toneR = `e;     15'd823: toneR = `e;
15'd824: toneR = `e;     15'd825: toneR = `e;
15'd826: toneR = `e;     15'd827: toneR = `e;
15'd828: toneR = `e;     15'd829: toneR = `e;
15'd830: toneR = `e;     15'd831: toneR = `e;
15'd832: toneR = `sil;     15'd833: toneR = `e;
15'd834: toneR = `e;     15'd835: toneR = `e;
15'd836: toneR = `f;     15'd837: toneR = `f;
15'd838: toneR = `f;     15'd839: toneR = `f;
15'd840: toneR = `g;     15'd841: toneR = `g;
15'd842: toneR = `g;     15'd843: toneR = `g;
15'd844: toneR = `g;     15'd845: toneR = `g;
15'd846: toneR = `g;     15'd847: toneR = `g;
15'd848: toneR = `sil;     15'd849: toneR = `g;
15'd850: toneR = `g;     15'd851: toneR = `g;
15'd852: toneR = `sil;     15'd853: toneR = `g;
15'd854: toneR = `g;     15'd855: toneR = `g;
15'd856: toneR = `g;     15'd857: toneR = `g;
15'd858: toneR = `g;     15'd859: toneR = `g;
15'd860: toneR = `sil;     15'd861: toneR = `g;
15'd862: toneR = `g;     15'd863: toneR = `g;
15'd864: toneR = `g;     15'd865: toneR = `g;
15'd866: toneR = `g;     15'd867: toneR = `g;
15'd868: toneR = `g;     15'd869: toneR = `g;
15'd870: toneR = `g;     15'd871: toneR = `g;
15'd872: toneR = `a;     15'd873: toneR = `a;
15'd874: toneR = `a;     15'd875: toneR = `a;
15'd876: toneR = `a;     15'd877: toneR = `a;
15'd878: toneR = `a;     15'd879: toneR = `a;
15'd880: toneR = `g;     15'd881: toneR = `g;
15'd882: toneR = `g;     15'd883: toneR = `g;
15'd884: toneR = `g;     15'd885: toneR = `g;
15'd886: toneR = `g;     15'd887: toneR = `g;
15'd888: toneR = `f;     15'd889: toneR = `f;
15'd890: toneR = `f;     15'd891: toneR = `f;
15'd892: toneR = `f;     15'd893: toneR = `f;
15'd894: toneR = `f;     15'd895: toneR = `f;
15'd896: toneR = `e;     15'd897: toneR = `e;
15'd898: toneR = `e;     15'd899: toneR = `e;
15'd900: toneR = `e;     15'd901: toneR = `e;
15'd902: toneR = `e;     15'd903: toneR = `e;
15'd904: toneR = `d;     15'd905: toneR = `d;
15'd906: toneR = `d;     15'd907: toneR = `d;
15'd908: toneR = `d;     15'd909: toneR = `d;
15'd910: toneR = `d;     15'd911: toneR = `d;
15'd912: toneR = `d;     15'd913: toneR = `d;
15'd914: toneR = `d;     15'd915: toneR = `d;
15'd916: toneR = `d;     15'd917: toneR = `d;
15'd918: toneR = `d;     15'd919: toneR = `d;
15'd920: toneR = `g;     15'd921: toneR = `g;
15'd922: toneR = `g;     15'd923: toneR = `g;
15'd924: toneR = `g;     15'd925: toneR = `g;
15'd926: toneR = `g;     15'd927: toneR = `g;
15'd928: toneR = `f;     15'd929: toneR = `f;
15'd930: toneR = `f;     15'd931: toneR = `f;
15'd932: toneR = `e;     15'd933: toneR = `e;
15'd934: toneR = `e;     15'd935: toneR = `e;
15'd936: toneR = `e;     15'd937: toneR = `e;
15'd938: toneR = `e;     15'd939: toneR = `e;
15'd940: toneR = `e;     15'd941: toneR = `e;
15'd942: toneR = `e;     15'd943: toneR = `e;
15'd944: toneR = `hc;     15'd945: toneR = `hc;
15'd946: toneR = `hc;     15'd947: toneR = `hc;
15'd948: toneR = `hc;     15'd949: toneR = `hc;
15'd950: toneR = `hc;     15'd951: toneR = `hc;
15'd952: toneR = `b;     15'd953: toneR = `b;
15'd954: toneR = `b;     15'd955: toneR = `b;
15'd956: toneR = `b;     15'd957: toneR = `b;
15'd958: toneR = `b;     15'd959: toneR = `b;
15'd960: toneR = `a;     15'd961: toneR = `a;
15'd962: toneR = `a;     15'd963: toneR = `a;
15'd964: toneR = `a;     15'd965: toneR = `a;
15'd966: toneR = `a;     15'd967: toneR = `a;
15'd968: toneR = `g;     15'd969: toneR = `g;
15'd970: toneR = `g;     15'd971: toneR = `g;
15'd972: toneR = `g;     15'd973: toneR = `g;
15'd974: toneR = `g;     15'd975: toneR = `g;
15'd976: toneR = `e;     15'd977: toneR = `e;
15'd978: toneR = `e;     15'd979: toneR = `e;
15'd980: toneR = `e;     15'd981: toneR = `e;
15'd982: toneR = `e;     15'd983: toneR = `e;
15'd984: toneR = `d;     15'd985: toneR = `d;
15'd986: toneR = `d;     15'd987: toneR = `d;
15'd988: toneR = `sil;     15'd989: toneR = `d;
15'd990: toneR = `d;     15'd991: toneR = `d;
15'd992: toneR = `d;     15'd993: toneR = `d;
15'd994: toneR = `d;     15'd995: toneR = `d;
15'd996: toneR = `d;     15'd997: toneR = `d;
15'd998: toneR = `d;     15'd999: toneR = `d;
15'd1000: toneR = `c;     15'd1001: toneR = `c;
15'd1002: toneR = `c;     15'd1003: toneR = `c;
15'd1004: toneR = `c;     15'd1005: toneR = `c;
15'd1006: toneR = `c;     15'd1007: toneR = `c;
15'd1008: toneR = `da;     15'd1009: toneR = `da;
15'd1010: toneR = `da;     15'd1011: toneR = `da;
15'd1012: toneR = `da;     15'd1013: toneR = `da;
15'd1014: toneR = `da;     15'd1015: toneR = `da;
15'd1016: toneR = `db;     15'd1017: toneR = `db;
15'd1018: toneR = `db;     15'd1019: toneR = `db;
15'd1020: toneR = `c;     15'd1021: toneR = `c;
15'd1022: toneR = `c;     15'd1023: toneR = `c;
15'd1024: toneR = `c;     15'd1025: toneR = `c;
15'd1026: toneR = `c;     15'd1027: toneR = `c;
15'd1028: toneR = `c;     15'd1029: toneR = `c;
15'd1030: toneR = `c;     15'd1031: toneR = `c;
15'd1032: toneR = `c;     15'd1033: toneR = `c;
15'd1034: toneR = `c;     15'd1035: toneR = `c;
15'd1036: toneR = `c;     15'd1037: toneR = `c;
15'd1038: toneR = `c;     15'd1039: toneR = `c;
15'd1040: toneR = `sil;     15'd1041: toneR = `sil;
15'd1042: toneR = `sil;     15'd1043: toneR = `sil;
15'd1044: toneR = `sil;     15'd1045: toneR = `sil;
15'd1046: toneR = `sil;     15'd1047: toneR = `sil;
15'd1048: toneR = `sil;     15'd1049: toneR = `sil;
15'd1050: toneR = `sil;     15'd1051: toneR = `sil;
15'd1052: toneR = `sil;     15'd1053: toneR = `sil;
15'd1054: toneR = `sil;     15'd1055: toneR = `sil;
15'd1056: toneR = `sil;     15'd1057: toneR = `sil;
15'd1058: toneR = `sil;     15'd1059: toneR = `sil;
15'd1060: toneR = `sil;     15'd1061: toneR = `sil;
15'd1062: toneR = `sil;     15'd1063: toneR = `sil;
15'd1064: toneR = `sil;     15'd1065: toneR = `sil;
15'd1066: toneR = `sil;     15'd1067: toneR = `sil;
15'd1068: toneR = `sil;     15'd1069: toneR = `sil;
15'd1070: toneR = `sil;     15'd1071: toneR = `sil;
15'd1072: toneR = `sil;     15'd1073: toneR = `sil;
15'd1074: toneR = `sil;     15'd1075: toneR = `sil;
15'd1076: toneR = `sil;     15'd1077: toneR = `sil;
15'd1078: toneR = `sil;     15'd1079: toneR = `sil;
15'd1080: toneR = `sil;     15'd1081: toneR = `sil;
15'd1082: toneR = `sil;     15'd1083: toneR = `sil;
15'd1084: toneR = `sil;     15'd1085: toneR = `sil;
15'd1086: toneR = `sil;     15'd1087: toneR = `sil;
15'd1088: toneR = `sil;     15'd1089: toneR = `sil;
15'd1090: toneR = `sil;     15'd1091: toneR = `sil;
15'd1092: toneR = `sil;     15'd1093: toneR = `sil;
15'd1094: toneR = `sil;     15'd1095: toneR = `sil;
15'd1096: toneR = `sil;     15'd1097: toneR = `sil;
15'd1098: toneR = `sil;     15'd1099: toneR = `sil;
15'd1100: toneR = `sil;     15'd1101: toneR = `sil;
15'd1102: toneR = `sil;     15'd1103: toneR = `sil;
15'd1104: toneR = `sil;     15'd1105: toneR = `sil;
15'd1106: toneR = `sil;     15'd1107: toneR = `sil;
15'd1108: toneR = `sil;     15'd1109: toneR = `sil;
15'd1110: toneR = `sil;     15'd1111: toneR = `sil;
15'd1112: toneR = `sil;     15'd1113: toneR = `sil;
15'd1114: toneR = `sil;     15'd1115: toneR = `sil;
15'd1116: toneR = `sil;     15'd1117: toneR = `sil;
15'd1118: toneR = `sil;     15'd1119: toneR = `sil;
15'd1120: toneR = `sil;     15'd1121: toneR = `sil;
15'd1122: toneR = `sil;     15'd1123: toneR = `sil;
15'd1124: toneR = `sil;     15'd1125: toneR = `sil;
15'd1126: toneR = `sil;     15'd1127: toneR = `sil;
15'd1128: toneR = `sil;     15'd1129: toneR = `sil;
15'd1130: toneR = `sil;     15'd1131: toneR = `sil;
15'd1132: toneR = `sil;     15'd1133: toneR = `sil;
15'd1134: toneR = `sil;     15'd1135: toneR = `sil;
15'd1136: toneR = `hc;     15'd1137: toneR = `hc;
15'd1138: toneR = `hc;     15'd1139: toneR = `hc;
15'd1140: toneR = `hc;     15'd1141: toneR = `hc;
15'd1142: toneR = `hc;     15'd1143: toneR = `hc;
15'd1144: toneR = `b;     15'd1145: toneR = `b;
15'd1146: toneR = `b;     15'd1147: toneR = `b;
15'd1148: toneR = `b;     15'd1149: toneR = `b;
15'd1150: toneR = `b;     15'd1151: toneR = `b;
15'd1152: toneR = `hc;     15'd1153: toneR = `hc;
15'd1154: toneR = `hc;     15'd1155: toneR = `hc;
15'd1156: toneR = `hc;     15'd1157: toneR = `hc;
15'd1158: toneR = `hc;     15'd1159: toneR = `hc;
15'd1160: toneR = `hc;     15'd1161: toneR = `hc;
15'd1162: toneR = `hc;     15'd1163: toneR = `hc;
15'd1164: toneR = `hc;     15'd1165: toneR = `hc;
15'd1166: toneR = `hc;     15'd1167: toneR = `hc;
15'd1168: toneR = `hc;     15'd1169: toneR = `hc;
15'd1170: toneR = `hc;     15'd1171: toneR = `hc;
15'd1172: toneR = `hc;     15'd1173: toneR = `hc;
15'd1174: toneR = `hc;     15'd1175: toneR = `hc;
15'd1176: toneR = `sil;     15'd1177: toneR = `hc;
15'd1178: toneR = `hc;     15'd1179: toneR = `hc;
15'd1180: toneR = `hc;     15'd1181: toneR = `hc;
15'd1182: toneR = `hc;     15'd1183: toneR = `hc;
15'd1184: toneR = `b;     15'd1185: toneR = `b;
15'd1186: toneR = `b;     15'd1187: toneR = `b;
15'd1188: toneR = `b;     15'd1189: toneR = `b;
15'd1190: toneR = `b;     15'd1191: toneR = `b;
15'd1192: toneR = `a;     15'd1193: toneR = `a;
15'd1194: toneR = `a;     15'd1195: toneR = `a;
15'd1196: toneR = `a;     15'd1197: toneR = `a;
15'd1198: toneR = `a;     15'd1199: toneR = `a;
15'd1200: toneR = `g;     15'd1201: toneR = `g;
15'd1202: toneR = `g;     15'd1203: toneR = `g;
15'd1204: toneR = `g;     15'd1205: toneR = `g;
15'd1206: toneR = `g;     15'd1207: toneR = `g;
15'd1208: toneR = `f;     15'd1209: toneR = `f;
15'd1210: toneR = `f;     15'd1211: toneR = `f;
15'd1212: toneR = `f;     15'd1213: toneR = `f;
15'd1214: toneR = `f;     15'd1215: toneR = `f;
                    default: toneR = `sil;
                endcase
            end
            else begin
                case(ibeatNum)
                    15'd0: toneR = `hc;     15'd1: toneR = `hc;
                    15'd2: toneR = `hc;     15'd3: toneR = `hc;
                    15'd4: toneR = `hc;     15'd5: toneR = `hc;
                    15'd6: toneR = `hc;     15'd7: toneR = `hc;
                    15'd8: toneR = `hc;     15'd9: toneR = `hc;
                    15'd10: toneR = `hc;     15'd11: toneR = `hc;
                    15'd12: toneR = `hc;     15'd13: toneR = `hc;
                    15'd14: toneR = `hc;     15'd15: toneR = `hc;
                    15'd16: toneR = `hd;     15'd17: toneR = `hd;
                    15'd18: toneR = `hd;     15'd19: toneR = `hd;
                    15'd20: toneR = `hd;     15'd21: toneR = `hd;
                    15'd22: toneR = `hd;     15'd23: toneR = `hd;
                    15'd24: toneR = `hd;     15'd25: toneR = `hd;
                    15'd26: toneR = `hd;     15'd27: toneR = `hd;
                    15'd28: toneR = `hd;     15'd29: toneR = `hd;
                    15'd30: toneR = `hd;     15'd31: toneR = `hd;
                    15'd32: toneR = `he;     15'd33: toneR = `he;
                    15'd34: toneR = `he;     15'd35: toneR = `he;
                    15'd36: toneR = `he;     15'd37: toneR = `he;
                    15'd38: toneR = `he;     15'd39: toneR = `he;
                    15'd40: toneR = `he;     15'd41: toneR = `he;
                    15'd42: toneR = `he;     15'd43: toneR = `he;
                    15'd44: toneR = `he;     15'd45: toneR = `he;
                    15'd46: toneR = `he;     15'd47: toneR = `he;
                    15'd48: toneR = `hc;     15'd49: toneR = `hc;
                    15'd50: toneR = `hc;     15'd51: toneR = `hc;
                    15'd52: toneR = `hc;     15'd53: toneR = `hc;
                    15'd54: toneR = `hc;     15'd55: toneR = `hc;
                    15'd56: toneR = `hc;     15'd57: toneR = `hc;
                    15'd58: toneR = `hc;     15'd59: toneR = `hc;
                    15'd60: toneR = `hc;     15'd61: toneR = `hc;
                    15'd62: toneR = `hc;     15'd63: toneR = `hc;
                    15'd64: toneR = `hc;     15'd65: toneR = `hc;
                    15'd66: toneR = `hc;     15'd67: toneR = `hc;
                    15'd68: toneR = `hc;     15'd69: toneR = `hc;
                    15'd70: toneR = `hc;     15'd71: toneR = `hc;
                    15'd72: toneR = `hc;     15'd73: toneR = `hc;
                    15'd74: toneR = `hc;     15'd75: toneR = `hc;
                    15'd76: toneR = `hc;     15'd77: toneR = `hc;
                    15'd78: toneR = `hc;     15'd79: toneR = `hc;
                    15'd80: toneR = `hd;     15'd81: toneR = `hd;
                    15'd82: toneR = `hd;     15'd83: toneR = `hd;
                    15'd84: toneR = `hd;     15'd85: toneR = `hd;
                    15'd86: toneR = `hd;     15'd87: toneR = `hd;
                    15'd88: toneR = `hd;     15'd89: toneR = `hd;
                    15'd90: toneR = `hd;     15'd91: toneR = `hd;
                    15'd92: toneR = `hd;     15'd93: toneR = `hd;
                    15'd94: toneR = `hd;     15'd95: toneR = `hd;
                    15'd96: toneR = `he;     15'd97: toneR = `he;
                    15'd98: toneR = `he;     15'd99: toneR = `he;
                    15'd100: toneR = `he;     15'd101: toneR = `he;
                    15'd102: toneR = `he;     15'd103: toneR = `he;
                    15'd104: toneR = `he;     15'd105: toneR = `he;
                    15'd106: toneR = `he;     15'd107: toneR = `he;
                    15'd108: toneR = `he;     15'd109: toneR = `he;
                    15'd110: toneR = `he;     15'd111: toneR = `he;
                    15'd112: toneR = `hc;     15'd113: toneR = `hc;
                    15'd114: toneR = `hc;     15'd115: toneR = `hc;
                    15'd116: toneR = `hc;     15'd117: toneR = `hc;
                    15'd118: toneR = `hc;     15'd119: toneR = `hc;
                    15'd120: toneR = `hc;     15'd121: toneR = `hc;
                    15'd122: toneR = `hc;     15'd123: toneR = `hc;
                    15'd124: toneR = `hc;     15'd125: toneR = `hc;
                    15'd126: toneR = `hc;     15'd127: toneR = `hc;
                    15'd128: toneR = `he;     15'd129: toneR = `he;
                    15'd130: toneR = `he;     15'd131: toneR = `he;
                    15'd132: toneR = `he;     15'd133: toneR = `he;
                    15'd134: toneR = `he;     15'd135: toneR = `he;
                    15'd136: toneR = `he;     15'd137: toneR = `he;
                    15'd138: toneR = `he;     15'd139: toneR = `he;
                    15'd140: toneR = `he;     15'd141: toneR = `he;
                    15'd142: toneR = `he;     15'd143: toneR = `he;
                    15'd144: toneR = `hf;     15'd145: toneR = `hf;
                    15'd146: toneR = `hf;     15'd147: toneR = `hf;
                    15'd148: toneR = `hf;     15'd149: toneR = `hf;
                    15'd150: toneR = `hf;     15'd151: toneR = `hf;
                    15'd152: toneR = `hf;     15'd153: toneR = `hf;
                    15'd154: toneR = `hf;     15'd155: toneR = `hf;
                    15'd156: toneR = `hf;     15'd157: toneR = `hf;
                    15'd158: toneR = `hf;     15'd159: toneR = `hf;
                    15'd160: toneR = `hg;     15'd161: toneR = `hg;
                    15'd162: toneR = `hg;     15'd163: toneR = `hg;
                    15'd164: toneR = `hg;     15'd165: toneR = `hg;
                    15'd166: toneR = `hg;     15'd167: toneR = `hg;
                    15'd168: toneR = `hg;     15'd169: toneR = `hg;
                    15'd170: toneR = `hg;     15'd171: toneR = `hg;
                    15'd172: toneR = `hg;     15'd173: toneR = `hg;
                    15'd174: toneR = `hg;     15'd175: toneR = `hg;
                    15'd176: toneR = `hg;     15'd177: toneR = `hg;
                    15'd178: toneR = `hg;     15'd179: toneR = `hg;
                    15'd180: toneR = `hg;     15'd181: toneR = `hg;
                    15'd182: toneR = `hg;     15'd183: toneR = `hg;
                    15'd184: toneR = `hg;     15'd185: toneR = `hg;
                    15'd186: toneR = `hg;     15'd187: toneR = `hg;
                    15'd188: toneR = `hg;     15'd189: toneR = `hg;
                    15'd190: toneR = `hg;     15'd191: toneR = `hg;
                    15'd192: toneR = `he;     15'd193: toneR = `he;
                    15'd194: toneR = `he;     15'd195: toneR = `he;
                    15'd196: toneR = `he;     15'd197: toneR = `he;
                    15'd198: toneR = `he;     15'd199: toneR = `he;
                    15'd200: toneR = `he;     15'd201: toneR = `he;
                    15'd202: toneR = `he;     15'd203: toneR = `he;
                    15'd204: toneR = `he;     15'd205: toneR = `he;
                    15'd206: toneR = `he;     15'd207: toneR = `he;
                    15'd208: toneR = `hf;     15'd209: toneR = `hf;
                    15'd210: toneR = `hf;     15'd211: toneR = `hf;
                    15'd212: toneR = `hf;     15'd213: toneR = `hf;
                    15'd214: toneR = `hf;     15'd215: toneR = `hf;
                    15'd216: toneR = `hf;     15'd217: toneR = `hf;
                    15'd218: toneR = `hf;     15'd219: toneR = `hf;
                    15'd220: toneR = `hf;     15'd221: toneR = `hf;
                    15'd222: toneR = `hf;     15'd223: toneR = `hf;
                    15'd224: toneR = `hg;     15'd225: toneR = `hg;
                    15'd226: toneR = `hg;     15'd227: toneR = `hg;
                    15'd228: toneR = `hg;     15'd229: toneR = `hg;
                    15'd230: toneR = `hg;     15'd231: toneR = `hg;
                    15'd232: toneR = `hg;     15'd233: toneR = `hg;
                    15'd234: toneR = `hg;     15'd235: toneR = `hg;
                    15'd236: toneR = `hg;     15'd237: toneR = `hg;
                    15'd238: toneR = `hg;     15'd239: toneR = `hg;
                    15'd240: toneR = `hg;     15'd241: toneR = `hg;
                    15'd242: toneR = `hg;     15'd243: toneR = `hg;
                    15'd244: toneR = `hg;     15'd245: toneR = `hg;
                    15'd246: toneR = `hg;     15'd247: toneR = `hg;
                    15'd248: toneR = `hg;     15'd249: toneR = `hg;
                    15'd250: toneR = `hg;     15'd251: toneR = `hg;
                    15'd252: toneR = `hg;     15'd253: toneR = `hg;
                    15'd254: toneR = `hg;     15'd255: toneR = `hg;
                    15'd256: toneR = `hg;     15'd257: toneR = `hg;
                    15'd258: toneR = `hg;     15'd259: toneR = `hg;
                    15'd260: toneR = `hg;     15'd261: toneR = `hg;
                    15'd262: toneR = `hg;     15'd263: toneR = `hg;
                    15'd264: toneR = `ha;     15'd265: toneR = `ha;
                    15'd266: toneR = `ha;     15'd267: toneR = `ha;
                    15'd268: toneR = `ha;     15'd269: toneR = `ha;
                    15'd270: toneR = `ha;     15'd271: toneR = `ha;
                    15'd272: toneR = `hg;     15'd273: toneR = `hg;
                    15'd274: toneR = `hg;     15'd275: toneR = `hg;
                    15'd276: toneR = `hg;     15'd277: toneR = `hg;
                    15'd278: toneR = `hg;     15'd279: toneR = `hg;
                    15'd280: toneR = `hf;     15'd281: toneR = `hf;
                    15'd282: toneR = `hf;     15'd283: toneR = `hf;
                    15'd284: toneR = `hf;     15'd285: toneR = `hf;
                    15'd286: toneR = `hf;     15'd287: toneR = `hf;
                    15'd288: toneR = `he;     15'd289: toneR = `he;
                    15'd290: toneR = `he;     15'd291: toneR = `he;
                    15'd292: toneR = `he;     15'd293: toneR = `he;
                    15'd294: toneR = `he;     15'd295: toneR = `he;
                    15'd296: toneR = `he;     15'd297: toneR = `he;
                    15'd298: toneR = `he;     15'd299: toneR = `he;
                    15'd300: toneR = `he;     15'd301: toneR = `he;
                    15'd302: toneR = `he;     15'd303: toneR = `he;
                    15'd304: toneR = `hc;     15'd305: toneR = `hc;
                    15'd306: toneR = `hc;     15'd307: toneR = `hc;
                    15'd308: toneR = `hc;     15'd309: toneR = `hc;
                    15'd310: toneR = `hc;     15'd311: toneR = `hc;
                    15'd312: toneR = `hc;     15'd313: toneR = `hc;
                    15'd314: toneR = `hc;     15'd315: toneR = `hc;
                    15'd316: toneR = `hc;     15'd317: toneR = `hc;
                    15'd318: toneR = `hc;     15'd319: toneR = `hc;
                    15'd320: toneR = `hg;     15'd321: toneR = `hg;
                    15'd322: toneR = `hg;     15'd323: toneR = `hg;
                    15'd324: toneR = `hg;     15'd325: toneR = `hg;
                    15'd326: toneR = `hg;     15'd327: toneR = `hg;
                    15'd328: toneR = `ha;     15'd329: toneR = `ha;
                    15'd330: toneR = `ha;     15'd331: toneR = `ha;
                    15'd332: toneR = `ha;     15'd333: toneR = `ha;
                    15'd334: toneR = `ha;     15'd335: toneR = `ha;
                    15'd336: toneR = `hg;     15'd337: toneR = `hg;
                    15'd338: toneR = `hg;     15'd339: toneR = `hg;
                    15'd340: toneR = `hg;     15'd341: toneR = `hg;
                    15'd342: toneR = `hg;     15'd343: toneR = `hg;
                    15'd344: toneR = `hf;     15'd345: toneR = `hf;
                    15'd346: toneR = `hf;     15'd347: toneR = `hf;
                    15'd348: toneR = `hf;     15'd349: toneR = `hf;
                    15'd350: toneR = `hf;     15'd351: toneR = `hf;
                    15'd352: toneR = `he;     15'd353: toneR = `he;
                    15'd354: toneR = `he;     15'd355: toneR = `he;
                    15'd356: toneR = `he;     15'd357: toneR = `he;
                    15'd358: toneR = `he;     15'd359: toneR = `he;
                    15'd360: toneR = `he;     15'd361: toneR = `he;
                    15'd362: toneR = `he;     15'd363: toneR = `he;
                    15'd364: toneR = `he;     15'd365: toneR = `he;
                    15'd366: toneR = `he;     15'd367: toneR = `he;
                    15'd368: toneR = `hc;     15'd369: toneR = `hc;
                    15'd370: toneR = `hc;     15'd371: toneR = `hc;
                    15'd372: toneR = `hc;     15'd373: toneR = `hc;
                    15'd374: toneR = `hc;     15'd375: toneR = `hc;
                    15'd376: toneR = `hc;     15'd377: toneR = `hc;
                    15'd378: toneR = `hc;     15'd379: toneR = `hc;
                    15'd380: toneR = `hc;     15'd381: toneR = `hc;
                    15'd382: toneR = `hc;     15'd383: toneR = `hc;
                    15'd384: toneR = `sil;     15'd385: toneR = `sil;
                    15'd386: toneR = `hc;     15'd387: toneR = `hc;
                    15'd388: toneR = `hc;     15'd389: toneR = `hc;
                    15'd390: toneR = `hc;     15'd391: toneR = `hc;
                    15'd392: toneR = `hc;     15'd393: toneR = `hc;
                    15'd394: toneR = `hc;     15'd395: toneR = `hc;
                    15'd396: toneR = `hc;     15'd397: toneR = `hc;
                    15'd398: toneR = `hc;     15'd399: toneR = `hc;
                    15'd400: toneR = `g;     15'd401: toneR = `g;
                    15'd402: toneR = `g;     15'd403: toneR = `g;
                    15'd404: toneR = `g;     15'd405: toneR = `g;
                    15'd406: toneR = `g;     15'd407: toneR = `g;
                    15'd408: toneR = `g;     15'd409: toneR = `g;
                    15'd410: toneR = `g;     15'd411: toneR = `g;
                    15'd412: toneR = `g;     15'd413: toneR = `g;
                    15'd414: toneR = `g;     15'd415: toneR = `g;
                    15'd416: toneR = `hc;     15'd417: toneR = `hc;
                    15'd418: toneR = `hc;     15'd419: toneR = `hc;
                    15'd420: toneR = `hc;     15'd421: toneR = `hc;
                    15'd422: toneR = `hc;     15'd423: toneR = `hc;
                    15'd424: toneR = `hc;     15'd425: toneR = `hc;
                    15'd426: toneR = `hc;     15'd427: toneR = `hc;
                    15'd428: toneR = `hc;     15'd429: toneR = `hc;
                    15'd430: toneR = `hc;     15'd431: toneR = `hc;
                    15'd432: toneR = `hc;     15'd433: toneR = `hc;
                    15'd434: toneR = `hc;     15'd435: toneR = `hc;
                    15'd436: toneR = `hc;     15'd437: toneR = `hc;
                    15'd438: toneR = `hc;     15'd439: toneR = `hc;
                    15'd440: toneR = `hc;     15'd441: toneR = `hc;
                    15'd442: toneR = `hc;     15'd443: toneR = `hc;
                    15'd444: toneR = `hc;     15'd445: toneR = `hc;
                    15'd446: toneR = `sil;     15'd447: toneR = `sil;
                    15'd448: toneR = `hc;     15'd449: toneR = `hc;
                    15'd450: toneR = `hc;     15'd451: toneR = `hc;
                    15'd452: toneR = `hc;     15'd453: toneR = `hc;
                    15'd454: toneR = `hc;     15'd455: toneR = `hc;
                    15'd456: toneR = `hc;     15'd457: toneR = `hc;
                    15'd458: toneR = `hc;     15'd459: toneR = `hc;
                    15'd460: toneR = `hc;     15'd461: toneR = `hc;
                    15'd462: toneR = `hc;     15'd463: toneR = `hc;
                    15'd464: toneR = `g;     15'd465: toneR = `g;
                    15'd466: toneR = `g;     15'd467: toneR = `g;
                    15'd468: toneR = `g;     15'd469: toneR = `g;
                    15'd470: toneR = `g;     15'd471: toneR = `g;
                    15'd472: toneR = `g;     15'd473: toneR = `g;
                    15'd474: toneR = `g;     15'd475: toneR = `g;
                    15'd476: toneR = `g;     15'd477: toneR = `g;
                    15'd478: toneR = `g;     15'd479: toneR = `g;
                    15'd480: toneR = `hc;     15'd481: toneR = `hc;
                    15'd482: toneR = `hc;     15'd483: toneR = `hc;
                    15'd484: toneR = `hc;     15'd485: toneR = `hc;
                    15'd486: toneR = `hc;     15'd487: toneR = `hc;
                    15'd488: toneR = `hc;     15'd489: toneR = `hc;
                    15'd490: toneR = `hc;     15'd491: toneR = `hc;
                    15'd492: toneR = `hc;     15'd493: toneR = `hc;
                    15'd494: toneR = `hc;     15'd495: toneR = `hc;
                    15'd496: toneR = `hc;     15'd497: toneR = `hc;
                    15'd498: toneR = `hc;     15'd499: toneR = `hc;
                    15'd500: toneR = `hc;     15'd501: toneR = `hc;
                    15'd502: toneR = `hc;     15'd503: toneR = `hc;
                    15'd504: toneR = `hc;     15'd505: toneR = `hc;
                    15'd506: toneR = `hc;     15'd507: toneR = `hc;
                    15'd508: toneR = `hc;     15'd509: toneR = `hc;
                    15'd510: toneR = `hc;     15'd511: toneR = `hc;
                    default: toneR = `sil;
                endcase
            end
            // case(ibeatNum)
                // // --- Measure 1 ---
                // 12'd0: toneR = `hg;      12'd1: toneR = `hg; // HG (half-beat)
                // 12'd2: toneR = `hg;      12'd3: toneR = `hg;
                // 12'd4: toneR = `hg;      12'd5: toneR = `hg;
                // 12'd6: toneR = `hg;      12'd7: toneR = `hg;
                // 12'd8: toneR = `he;      12'd9: toneR = `he; // HE (half-beat)
                // 12'd10: toneR = `he;     12'd11: toneR = `he;
                // 12'd12: toneR = `he;     12'd13: toneR = `he;
                // 12'd14: toneR = `he;     12'd15: toneR = `sil; // (Short break for repetitive notes: high E)

                // 12'd16: toneR = `he;     12'd17: toneR = `he; // HE (one-beat)
                // 12'd18: toneR = `he;     12'd19: toneR = `he;
                // 12'd20: toneR = `he;     12'd21: toneR = `he;
                // 12'd22: toneR = `he;     12'd23: toneR = `he;
                // 12'd24: toneR = `he;     12'd25: toneR = `he;
                // 12'd26: toneR = `he;     12'd27: toneR = `he;
                // 12'd28: toneR = `he;     12'd29: toneR = `he;
                // 12'd30: toneR = `he;     12'd31: toneR = `he;

                // 12'd32: toneR = `hf;     12'd33: toneR = `hf; // HF (half-beat)
                // 12'd34: toneR = `hf;     12'd35: toneR = `hf;
                // 12'd36: toneR = `hf;     12'd37: toneR = `hf;
                // 12'd38: toneR = `hf;     12'd39: toneR = `hf;
                // 12'd40: toneR = `hd;     12'd41: toneR = `hd; // HD (half-beat)
                // 12'd42: toneR = `hd;     12'd43: toneR = `hd;
                // 12'd44: toneR = `hd;     12'd45: toneR = `hd;
                // 12'd46: toneR = `hd;     12'd47: toneR = `sil; // (Short break for repetitive notes: high D)

                // 12'd48: toneR = `hd;     12'd49: toneR = `hd; // HD (one-beat)
                // 12'd50: toneR = `hd;     12'd51: toneR = `hd;
                // 12'd52: toneR = `hd;     12'd53: toneR = `hd;
                // 12'd54: toneR = `hd;     12'd55: toneR = `hd;
                // 12'd56: toneR = `hd;     12'd57: toneR = `hd;
                // 12'd58: toneR = `hd;     12'd59: toneR = `hd;
                // 12'd60: toneR = `hd;     12'd61: toneR = `hd;
                // 12'd62: toneR = `hd;     12'd63: toneR = `hd;

                // // --- Measure 2 ---
                // 12'd64: toneR = `hc;     12'd65: toneR = `hc; // HC (half-beat)
                // 12'd66: toneR = `hc;     12'd67: toneR = `hc;
                // 12'd68: toneR = `hc;     12'd69: toneR = `hc;
                // 12'd70: toneR = `hc;     12'd71: toneR = `hc;
                // 12'd72: toneR = `hd;     12'd73: toneR = `hd; // HD (half-beat)
                // 12'd74: toneR = `hd;     12'd75: toneR = `hd;
                // 12'd76: toneR = `hd;     12'd77: toneR = `hd;
                // 12'd78: toneR = `hd;     12'd79: toneR = `hd;

                // 12'd80: toneR = `he;     12'd81: toneR = `he; // HE (half-beat)
                // 12'd82: toneR = `he;     12'd83: toneR = `he;
                // 12'd84: toneR = `he;     12'd85: toneR = `he;
                // 12'd86: toneR = `he;     12'd87: toneR = `he;
                // 12'd88: toneR = `hf;     12'd89: toneR = `hf; // HF (half-beat)
                // 12'd90: toneR = `hf;     12'd91: toneR = `hf;
                // 12'd92: toneR = `hf;     12'd93: toneR = `hf;
                // 12'd94: toneR = `hf;     12'd95: toneR = `hf;

                // 12'd96: toneR = `hg;     12'd97: toneR = `hg; // HG (half-beat)
                // 12'd98: toneR = `hg;     12'd99: toneR = `hg;
                // 12'd100: toneR = `hg;     12'd101: toneR = `hg;
                // 12'd102: toneR = `hg;     12'd103: toneR = `sil; // (Short break for repetitive notes: high D)
                // 12'd104: toneR = `hg;     12'd105: toneR = `hg; // HG (half-beat)
                // 12'd106: toneR = `hg;     12'd107: toneR = `hg;
                // 12'd108: toneR = `hg;     12'd109: toneR = `hg;
                // 12'd110: toneR = `hg;     12'd111: toneR = `sil; // (Short break for repetitive notes: high D)

                // 12'd112: toneR = `hg;     12'd113: toneR = `hg; // HG (one-beat)
                // 12'd114: toneR = `hg;     12'd115: toneR = `hg;
                // 12'd116: toneR = `hg;     12'd117: toneR = `hg;
                // 12'd118: toneR = `hg;     12'd119: toneR = `hg;
                // 12'd120: toneR = `hg;     12'd121: toneR = `hg;
                // 12'd122: toneR = `hg;     12'd123: toneR = `hg;
                // 12'd124: toneR = `hg;     12'd125: toneR = `hg;
                // 12'd126: toneR = `hg;     12'd127: toneR = `hg;

                // 15'd0: toneR = `ha;     15'd1: toneR = `ha;
                // 15'd2: toneR = `ha;     15'd3: toneR = `ha;
                // 15'd4: toneR = `ha;     15'd5: toneR = `ha;
                // 15'd6: toneR = `ha;     15'd7: toneR = `ha;
                // 15'd8: toneR = `rhf;     15'd9: toneR = `rhf;
                // 15'd10: toneR = `rhf;     15'd11: toneR = `rhf;
                // 15'd12: toneR = `hg;     15'd13: toneR = `hg;
                // 15'd14: toneR = `hg;     15'd15: toneR = `hg;
                // 15'd16: toneR = `ha;     15'd17: toneR = `ha;
                // 15'd18: toneR = `ha;     15'd19: toneR = `ha;
                // 15'd20: toneR = `ha;     15'd21: toneR = `ha;
                // 15'd22: toneR = `ha;     15'd23: toneR = `ha;
                // 15'd24: toneR = `rhf;     15'd25: toneR = `rhf;
                // 15'd26: toneR = `rhf;     15'd27: toneR = `rhf;
                // 15'd28: toneR = `hg;     15'd29: toneR = `hg;
                // 15'd30: toneR = `hg;     15'd31: toneR = `hg;
                // 15'd32: toneR = `ha;     15'd33: toneR = `ha;
                // 15'd34: toneR = `ha;     15'd35: toneR = `ha;
                // 15'd36: toneR = `a;     15'd37: toneR = `a;
                // 15'd38: toneR = `a;     15'd39: toneR = `a;
                // 15'd40: toneR = `b;     15'd41: toneR = `b;
                // 15'd42: toneR = `b;     15'd43: toneR = `b;
                // 15'd44: toneR = `rhc;     15'd45: toneR = `rhc;
                // 15'd46: toneR = `rhc;     15'd47: toneR = `rhc;
                // 15'd48: toneR = `hd;     15'd49: toneR = `hd;
                // 15'd50: toneR = `hd;     15'd51: toneR = `hd;
                // 15'd52: toneR = `he;     15'd53: toneR = `he;
                // 15'd54: toneR = `he;     15'd55: toneR = `he;
                // 15'd56: toneR = `rhf;     15'd57: toneR = `rhf;
                // 15'd58: toneR = `rhf;     15'd59: toneR = `rhf;
                // 15'd60: toneR = `hg;     15'd61: toneR = `hg;
                // 15'd62: toneR = `hg;     15'd63: toneR = `hg;
                // 15'd64: toneR = `rhf;     15'd65: toneR = `rhf;
                // 15'd66: toneR = `rhf;     15'd67: toneR = `rhf;
                // 15'd68: toneR = `rhf;     15'd69: toneR = `rhf;
                // 15'd70: toneR = `rhf;     15'd71: toneR = `rhf;
                // 15'd72: toneR = `hd;     15'd73: toneR = `hd;
                // 15'd74: toneR = `hd;     15'd75: toneR = `hd;
                // 15'd76: toneR = `he;     15'd77: toneR = `he;
                // 15'd78: toneR = `he;     15'd79: toneR = `he;
                // 15'd80: toneR = `rhf;     15'd81: toneR = `rhf;
                // 15'd82: toneR = `rhf;     15'd83: toneR = `rhf;
                // 15'd84: toneR = `rhf;     15'd85: toneR = `rhf;
                // 15'd86: toneR = `rhf;     15'd87: toneR = `rhf;
                // 15'd88: toneR = `rf;     15'd89: toneR = `rf;
                // 15'd90: toneR = `rf;     15'd91: toneR = `rf;
                // 15'd92: toneR = `g;     15'd93: toneR = `g;
                // 15'd94: toneR = `g;     15'd95: toneR = `g;
                // 15'd96: toneR = `a;     15'd97: toneR = `a;
                // 15'd98: toneR = `a;     15'd99: toneR = `a;
                // 15'd100: toneR = `b;     15'd101: toneR = `b;
                // 15'd102: toneR = `b;     15'd103: toneR = `b;
                // 15'd104: toneR = `a;     15'd105: toneR = `a;
                // 15'd106: toneR = `a;     15'd107: toneR = `a;
                // 15'd108: toneR = `g;     15'd109: toneR = `g;
                // 15'd110: toneR = `g;     15'd111: toneR = `g;
                // 15'd112: toneR = `a;     15'd113: toneR = `a;
                // 15'd114: toneR = `a;     15'd115: toneR = `a;
                // 15'd116: toneR = `rf;     15'd117: toneR = `rf;
                // 15'd118: toneR = `rf;     15'd119: toneR = `rf;
                // 15'd120: toneR = `g;     15'd121: toneR = `g;
                // 15'd122: toneR = `g;     15'd123: toneR = `g;
                // 15'd124: toneR = `a;     15'd125: toneR = `a;
                // 15'd126: toneR = `a;     15'd127: toneR = `a;
                // 15'd128: toneR = `g;     15'd129: toneR = `g;
                // 15'd130: toneR = `g;     15'd131: toneR = `g;
                // 15'd132: toneR = `g;     15'd133: toneR = `g;
                // 15'd134: toneR = `g;     15'd135: toneR = `g;
                // 15'd136: toneR = `b;     15'd137: toneR = `b;
                // 15'd138: toneR = `b;     15'd139: toneR = `b;
                // 15'd140: toneR = `a;     15'd141: toneR = `a;
                // 15'd142: toneR = `a;     15'd143: toneR = `a;
                // 15'd144: toneR = `g;     15'd145: toneR = `g;
                // 15'd146: toneR = `g;     15'd147: toneR = `g;
                // 15'd148: toneR = `g;     15'd149: toneR = `g;
                // 15'd150: toneR = `g;     15'd151: toneR = `g;
                // 15'd152: toneR = `rf;     15'd153: toneR = `rf;
                // 15'd154: toneR = `rf;     15'd155: toneR = `rf;
                // 15'd156: toneR = `e;     15'd157: toneR = `e;
                // 15'd158: toneR = `e;     15'd159: toneR = `e;
                // 15'd160: toneR = `rf;     15'd161: toneR = `rf;
                // 15'd162: toneR = `rf;     15'd163: toneR = `rf;
                // 15'd164: toneR = `e;     15'd165: toneR = `e;
                // 15'd166: toneR = `e;     15'd167: toneR = `e;
                // 15'd168: toneR = `d;     15'd169: toneR = `d;
                // 15'd170: toneR = `d;     15'd171: toneR = `d;
                // 15'd172: toneR = `e;     15'd173: toneR = `e;
                // 15'd174: toneR = `e;     15'd175: toneR = `e;
                // 15'd176: toneR = `rf;     15'd177: toneR = `rf;
                // 15'd178: toneR = `rf;     15'd179: toneR = `rf;
                // 15'd180: toneR = `g;     15'd181: toneR = `g;
                // 15'd182: toneR = `g;     15'd183: toneR = `g;
                // 15'd184: toneR = `a;     15'd185: toneR = `a;
                // 15'd186: toneR = `a;     15'd187: toneR = `a;
                // 15'd188: toneR = `b;     15'd189: toneR = `b;
                // 15'd190: toneR = `b;     15'd191: toneR = `b;
                // 15'd192: toneR = `g;     15'd193: toneR = `g;
                // 15'd194: toneR = `g;     15'd195: toneR = `g;
                // 15'd196: toneR = `g;     15'd197: toneR = `g;
                // 15'd198: toneR = `g;     15'd199: toneR = `g;
                // 15'd200: toneR = `b;     15'd201: toneR = `b;
                // 15'd202: toneR = `b;     15'd203: toneR = `b;
                // 15'd204: toneR = `a;     15'd205: toneR = `a;
                // 15'd206: toneR = `a;     15'd207: toneR = `a;
                // 15'd208: toneR = `b;     15'd209: toneR = `b;
                // 15'd210: toneR = `b;     15'd211: toneR = `b;
                // 15'd212: toneR = `b;     15'd213: toneR = `b;
                // 15'd214: toneR = `b;     15'd215: toneR = `b;
                // 15'd216: toneR = `rhc;     15'd217: toneR = `rhc;
                // 15'd218: toneR = `rhc;     15'd219: toneR = `rhc;
                // 15'd220: toneR = `hd;     15'd221: toneR = `hd;
                // 15'd222: toneR = `hd;     15'd223: toneR = `hd;
                // 15'd224: toneR = `a;     15'd225: toneR = `a;
                // 15'd226: toneR = `a;     15'd227: toneR = `a;
                // 15'd228: toneR = `b;     15'd229: toneR = `b;
                // 15'd230: toneR = `b;     15'd231: toneR = `b;
                // 15'd232: toneR = `rhc;     15'd233: toneR = `rhc;
                // 15'd234: toneR = `rhc;     15'd235: toneR = `rhc;
                // 15'd236: toneR = `hd;     15'd237: toneR = `hd;
                // 15'd238: toneR = `hd;     15'd239: toneR = `hd;
                // 15'd240: toneR = `he;     15'd241: toneR = `he;
                // 15'd242: toneR = `he;     15'd243: toneR = `he;
                // 15'd244: toneR = `rhf;     15'd245: toneR = `rhf;
                // 15'd246: toneR = `rhf;     15'd247: toneR = `rhf;
                // 15'd248: toneR = `hg;     15'd249: toneR = `hg;
                // 15'd250: toneR = `hg;     15'd251: toneR = `hg;
                // 15'd252: toneR = `ha;     15'd253: toneR = `ha;
                // 15'd254: toneR = `ha;     15'd255: toneR = `ha;
                // 15'd256: toneR = `rhf;     15'd257: toneR = `rhf;
                // 15'd258: toneR = `rhf;     15'd259: toneR = `rhf;
                // 15'd260: toneR = `rhf;     15'd261: toneR = `rhf;
                // 15'd262: toneR = `rhf;     15'd263: toneR = `rhf;
                // 15'd264: toneR = `hd;     15'd265: toneR = `hd;
                // 15'd266: toneR = `hd;     15'd267: toneR = `hd;
                // 15'd268: toneR = `he;     15'd269: toneR = `he;
                // 15'd270: toneR = `he;     15'd271: toneR = `he;
                // 15'd272: toneR = `rhf;     15'd273: toneR = `rhf;
                // 15'd274: toneR = `rhf;     15'd275: toneR = `rhf;
                // 15'd276: toneR = `rhf;     15'd277: toneR = `rhf;
                // 15'd278: toneR = `rhf;     15'd279: toneR = `rhf;
                // 15'd280: toneR = `he;     15'd281: toneR = `he;
                // 15'd282: toneR = `he;     15'd283: toneR = `he;
                // 15'd284: toneR = `hd;     15'd285: toneR = `hd;
                // 15'd286: toneR = `hd;     15'd287: toneR = `hd;
                // 15'd288: toneR = `he;     15'd289: toneR = `he;
                // 15'd290: toneR = `he;     15'd291: toneR = `he;
                // 15'd292: toneR = `rhc;     15'd293: toneR = `rhc;
                // 15'd294: toneR = `rhc;     15'd295: toneR = `rhc;
                // 15'd296: toneR = `hd;     15'd297: toneR = `hd;
                // 15'd298: toneR = `hd;     15'd299: toneR = `hd;
                // 15'd300: toneR = `he;     15'd301: toneR = `he;
                // 15'd302: toneR = `he;     15'd303: toneR = `he;
                // 15'd304: toneR = `rhf;     15'd305: toneR = `rhf;
                // 15'd306: toneR = `rhf;     15'd307: toneR = `rhf;
                // 15'd308: toneR = `he;     15'd309: toneR = `he;
                // 15'd310: toneR = `he;     15'd311: toneR = `he;
                // 15'd312: toneR = `hd;     15'd313: toneR = `hd;
                // 15'd314: toneR = `hd;     15'd315: toneR = `hd;
                // 15'd316: toneR = `rhc;     15'd317: toneR = `rhc;
                // 15'd318: toneR = `rhc;     15'd319: toneR = `rhc;

        //         15'd0: toneR = `hc;     15'd1: toneR = `hc;
        //             15'd2: toneR = `hc;     15'd3: toneR = `hc;
        //             15'd4: toneR = `hc;     15'd5: toneR = `hc;
        //             15'd6: toneR = `hc;     15'd7: toneR = `hc;
        //             15'd8: toneR = `hc;     15'd9: toneR = `hc;
        //             15'd10: toneR = `hc;     15'd11: toneR = `hc;
        //             15'd12: toneR = `hc;     15'd13: toneR = `hc;
        //             15'd14: toneR = `hc;     15'd15: toneR = `hc;
        //             15'd16: toneR = `hd;     15'd17: toneR = `hd;
        //             15'd18: toneR = `hd;     15'd19: toneR = `hd;
        //             15'd20: toneR = `hd;     15'd21: toneR = `hd;
        //             15'd22: toneR = `hd;     15'd23: toneR = `hd;
        //             15'd24: toneR = `hd;     15'd25: toneR = `hd;
        //             15'd26: toneR = `hd;     15'd27: toneR = `hd;
        //             15'd28: toneR = `hd;     15'd29: toneR = `hd;
        //             15'd30: toneR = `hd;     15'd31: toneR = `hd;
        //             15'd32: toneR = `he;     15'd33: toneR = `he;
        //             15'd34: toneR = `he;     15'd35: toneR = `he;
        //             15'd36: toneR = `he;     15'd37: toneR = `he;
        //             15'd38: toneR = `he;     15'd39: toneR = `he;
        //             15'd40: toneR = `he;     15'd41: toneR = `he;
        //             15'd42: toneR = `he;     15'd43: toneR = `he;
        //             15'd44: toneR = `he;     15'd45: toneR = `he;
        //             15'd46: toneR = `he;     15'd47: toneR = `he;
        //             15'd48: toneR = `hc;     15'd49: toneR = `hc;
        //             15'd50: toneR = `hc;     15'd51: toneR = `hc;
        //             15'd52: toneR = `hc;     15'd53: toneR = `hc;
        //             15'd54: toneR = `hc;     15'd55: toneR = `hc;
        //             15'd56: toneR = `hc;     15'd57: toneR = `hc;
        //             15'd58: toneR = `hc;     15'd59: toneR = `hc;
        //             15'd60: toneR = `hc;     15'd61: toneR = `hc;
        //             15'd62: toneR = `hc;     15'd63: toneR = `hc;
        //             15'd64: toneR = `hc;     15'd65: toneR = `hc;
        //             15'd66: toneR = `hc;     15'd67: toneR = `hc;
        //             15'd68: toneR = `hc;     15'd69: toneR = `hc;
        //             15'd70: toneR = `hc;     15'd71: toneR = `hc;
        //             15'd72: toneR = `hc;     15'd73: toneR = `hc;
        //             15'd74: toneR = `hc;     15'd75: toneR = `hc;
        //             15'd76: toneR = `hc;     15'd77: toneR = `hc;
        //             15'd78: toneR = `hc;     15'd79: toneR = `hc;
        //             15'd80: toneR = `hd;     15'd81: toneR = `hd;
        //             15'd82: toneR = `hd;     15'd83: toneR = `hd;
        //             15'd84: toneR = `hd;     15'd85: toneR = `hd;
        //             15'd86: toneR = `hd;     15'd87: toneR = `hd;
        //             15'd88: toneR = `hd;     15'd89: toneR = `hd;
        //             15'd90: toneR = `hd;     15'd91: toneR = `hd;
        //             15'd92: toneR = `hd;     15'd93: toneR = `hd;
        //             15'd94: toneR = `hd;     15'd95: toneR = `hd;
        //             15'd96: toneR = `he;     15'd97: toneR = `he;
        //             15'd98: toneR = `he;     15'd99: toneR = `he;
        //             15'd100: toneR = `he;     15'd101: toneR = `he;
        //             15'd102: toneR = `he;     15'd103: toneR = `he;
        //             15'd104: toneR = `he;     15'd105: toneR = `he;
        //             15'd106: toneR = `he;     15'd107: toneR = `he;
        //             15'd108: toneR = `he;     15'd109: toneR = `he;
        //             15'd110: toneR = `he;     15'd111: toneR = `he;
        //             15'd112: toneR = `hc;     15'd113: toneR = `hc;
        //             15'd114: toneR = `hc;     15'd115: toneR = `hc;
        //             15'd116: toneR = `hc;     15'd117: toneR = `hc;
        //             15'd118: toneR = `hc;     15'd119: toneR = `hc;
        //             15'd120: toneR = `hc;     15'd121: toneR = `hc;
        //             15'd122: toneR = `hc;     15'd123: toneR = `hc;
        //             15'd124: toneR = `hc;     15'd125: toneR = `hc;
        //             15'd126: toneR = `hc;     15'd127: toneR = `hc;
        //             15'd128: toneR = `he;     15'd129: toneR = `he;
        //             15'd130: toneR = `he;     15'd131: toneR = `he;
        //             15'd132: toneR = `he;     15'd133: toneR = `he;
        //             15'd134: toneR = `he;     15'd135: toneR = `he;
        //             15'd136: toneR = `he;     15'd137: toneR = `he;
        //             15'd138: toneR = `he;     15'd139: toneR = `he;
        //             15'd140: toneR = `he;     15'd141: toneR = `he;
        //             15'd142: toneR = `he;     15'd143: toneR = `he;
        //             15'd144: toneR = `hf;     15'd145: toneR = `hf;
        //             15'd146: toneR = `hf;     15'd147: toneR = `hf;
        //             15'd148: toneR = `hf;     15'd149: toneR = `hf;
        //             15'd150: toneR = `hf;     15'd151: toneR = `hf;
        //             15'd152: toneR = `hf;     15'd153: toneR = `hf;
        //             15'd154: toneR = `hf;     15'd155: toneR = `hf;
        //             15'd156: toneR = `hf;     15'd157: toneR = `hf;
        //             15'd158: toneR = `hf;     15'd159: toneR = `hf;
        //             15'd160: toneR = `hg;     15'd161: toneR = `hg;
        //             15'd162: toneR = `hg;     15'd163: toneR = `hg;
        //             15'd164: toneR = `hg;     15'd165: toneR = `hg;
        //             15'd166: toneR = `hg;     15'd167: toneR = `hg;
        //             15'd168: toneR = `hg;     15'd169: toneR = `hg;
        //             15'd170: toneR = `hg;     15'd171: toneR = `hg;
        //             15'd172: toneR = `hg;     15'd173: toneR = `hg;
        //             15'd174: toneR = `hg;     15'd175: toneR = `hg;
        //             15'd176: toneR = `hg;     15'd177: toneR = `hg;
        //             15'd178: toneR = `hg;     15'd179: toneR = `hg;
        //             15'd180: toneR = `hg;     15'd181: toneR = `hg;
        //             15'd182: toneR = `hg;     15'd183: toneR = `hg;
        //             15'd184: toneR = `hg;     15'd185: toneR = `hg;
        //             15'd186: toneR = `hg;     15'd187: toneR = `hg;
        //             15'd188: toneR = `hg;     15'd189: toneR = `hg;
        //             15'd190: toneR = `hg;     15'd191: toneR = `hg;
        //             15'd192: toneR = `he;     15'd193: toneR = `he;
        //             15'd194: toneR = `he;     15'd195: toneR = `he;
        //             15'd196: toneR = `he;     15'd197: toneR = `he;
        //             15'd198: toneR = `he;     15'd199: toneR = `he;
        //             15'd200: toneR = `he;     15'd201: toneR = `he;
        //             15'd202: toneR = `he;     15'd203: toneR = `he;
        //             15'd204: toneR = `he;     15'd205: toneR = `he;
        //             15'd206: toneR = `he;     15'd207: toneR = `he;
        //             15'd208: toneR = `hf;     15'd209: toneR = `hf;
        //             15'd210: toneR = `hf;     15'd211: toneR = `hf;
        //             15'd212: toneR = `hf;     15'd213: toneR = `hf;
        //             15'd214: toneR = `hf;     15'd215: toneR = `hf;
        //             15'd216: toneR = `hf;     15'd217: toneR = `hf;
        //             15'd218: toneR = `hf;     15'd219: toneR = `hf;
        //             15'd220: toneR = `hf;     15'd221: toneR = `hf;
        //             15'd222: toneR = `hf;     15'd223: toneR = `hf;
        //             15'd224: toneR = `hg;     15'd225: toneR = `hg;
        //             15'd226: toneR = `hg;     15'd227: toneR = `hg;
        //             15'd228: toneR = `hg;     15'd229: toneR = `hg;
        //             15'd230: toneR = `hg;     15'd231: toneR = `hg;
        //             15'd232: toneR = `hg;     15'd233: toneR = `hg;
        //             15'd234: toneR = `hg;     15'd235: toneR = `hg;
        //             15'd236: toneR = `hg;     15'd237: toneR = `hg;
        //             15'd238: toneR = `hg;     15'd239: toneR = `hg;
        //             15'd240: toneR = `hg;     15'd241: toneR = `hg;
        //             15'd242: toneR = `hg;     15'd243: toneR = `hg;
        //             15'd244: toneR = `hg;     15'd245: toneR = `hg;
        //             15'd246: toneR = `hg;     15'd247: toneR = `hg;
        //             15'd248: toneR = `hg;     15'd249: toneR = `hg;
        //             15'd250: toneR = `hg;     15'd251: toneR = `hg;
        //             15'd252: toneR = `hg;     15'd253: toneR = `hg;
        //             15'd254: toneR = `hg;     15'd255: toneR = `hg;
        //             15'd256: toneR = `hg;     15'd257: toneR = `hg;
        //             15'd258: toneR = `hg;     15'd259: toneR = `hg;
        //             15'd260: toneR = `hg;     15'd261: toneR = `hg;
        //             15'd262: toneR = `hg;     15'd263: toneR = `hg;
        //             15'd264: toneR = `ha;     15'd265: toneR = `ha;
        //             15'd266: toneR = `ha;     15'd267: toneR = `ha;
        //             15'd268: toneR = `ha;     15'd269: toneR = `ha;
        //             15'd270: toneR = `ha;     15'd271: toneR = `ha;
        //             15'd272: toneR = `hg;     15'd273: toneR = `hg;
        //             15'd274: toneR = `hg;     15'd275: toneR = `hg;
        //             15'd276: toneR = `hg;     15'd277: toneR = `hg;
        //             15'd278: toneR = `hg;     15'd279: toneR = `hg;
        //             15'd280: toneR = `hf;     15'd281: toneR = `hf;
        //             15'd282: toneR = `hf;     15'd283: toneR = `hf;
        //             15'd284: toneR = `hf;     15'd285: toneR = `hf;
        //             15'd286: toneR = `hf;     15'd287: toneR = `hf;
        //             15'd288: toneR = `he;     15'd289: toneR = `he;
        //             15'd290: toneR = `he;     15'd291: toneR = `he;
        //             15'd292: toneR = `he;     15'd293: toneR = `he;
        //             15'd294: toneR = `he;     15'd295: toneR = `he;
        //             15'd296: toneR = `he;     15'd297: toneR = `he;
        //             15'd298: toneR = `he;     15'd299: toneR = `he;
        //             15'd300: toneR = `he;     15'd301: toneR = `he;
        //             15'd302: toneR = `he;     15'd303: toneR = `he;
        //             15'd304: toneR = `hc;     15'd305: toneR = `hc;
        //             15'd306: toneR = `hc;     15'd307: toneR = `hc;
        //             15'd308: toneR = `hc;     15'd309: toneR = `hc;
        //             15'd310: toneR = `hc;     15'd311: toneR = `hc;
        //             15'd312: toneR = `hc;     15'd313: toneR = `hc;
        //             15'd314: toneR = `hc;     15'd315: toneR = `hc;
        //             15'd316: toneR = `hc;     15'd317: toneR = `hc;
        //             15'd318: toneR = `hc;     15'd319: toneR = `hc;
        //             15'd320: toneR = `hg;     15'd321: toneR = `hg;
        //             15'd322: toneR = `hg;     15'd323: toneR = `hg;
        //             15'd324: toneR = `hg;     15'd325: toneR = `hg;
        //             15'd326: toneR = `hg;     15'd327: toneR = `hg;
        //             15'd328: toneR = `ha;     15'd329: toneR = `ha;
        //             15'd330: toneR = `ha;     15'd331: toneR = `ha;
        //             15'd332: toneR = `ha;     15'd333: toneR = `ha;
        //             15'd334: toneR = `ha;     15'd335: toneR = `ha;
        //             15'd336: toneR = `hg;     15'd337: toneR = `hg;
        //             15'd338: toneR = `hg;     15'd339: toneR = `hg;
        //             15'd340: toneR = `hg;     15'd341: toneR = `hg;
        //             15'd342: toneR = `hg;     15'd343: toneR = `hg;
        //             15'd344: toneR = `hf;     15'd345: toneR = `hf;
        //             15'd346: toneR = `hf;     15'd347: toneR = `hf;
        //             15'd348: toneR = `hf;     15'd349: toneR = `hf;
        //             15'd350: toneR = `hf;     15'd351: toneR = `hf;
        //             15'd352: toneR = `he;     15'd353: toneR = `he;
        //             15'd354: toneR = `he;     15'd355: toneR = `he;
        //             15'd356: toneR = `he;     15'd357: toneR = `he;
        //             15'd358: toneR = `he;     15'd359: toneR = `he;
        //             15'd360: toneR = `he;     15'd361: toneR = `he;
        //             15'd362: toneR = `he;     15'd363: toneR = `he;
        //             15'd364: toneR = `he;     15'd365: toneR = `he;
        //             15'd366: toneR = `he;     15'd367: toneR = `he;
        //             15'd368: toneR = `hc;     15'd369: toneR = `hc;
        //             15'd370: toneR = `hc;     15'd371: toneR = `hc;
        //             15'd372: toneR = `hc;     15'd373: toneR = `hc;
        //             15'd374: toneR = `hc;     15'd375: toneR = `hc;
        //             15'd376: toneR = `hc;     15'd377: toneR = `hc;
        //             15'd378: toneR = `hc;     15'd379: toneR = `hc;
        //             15'd380: toneR = `hc;     15'd381: toneR = `hc;
        //             15'd382: toneR = `hc;     15'd383: toneR = `hc;
        //             15'd384: toneR = `sil;     15'd385: toneR = `sil;
        //             15'd386: toneR = `hc;     15'd387: toneR = `hc;
        //             15'd388: toneR = `hc;     15'd389: toneR = `hc;
        //             15'd390: toneR = `hc;     15'd391: toneR = `hc;
        //             15'd392: toneR = `hc;     15'd393: toneR = `hc;
        //             15'd394: toneR = `hc;     15'd395: toneR = `hc;
        //             15'd396: toneR = `hc;     15'd397: toneR = `hc;
        //             15'd398: toneR = `hc;     15'd399: toneR = `hc;
        //             15'd400: toneR = `g;     15'd401: toneR = `g;
        //             15'd402: toneR = `g;     15'd403: toneR = `g;
        //             15'd404: toneR = `g;     15'd405: toneR = `g;
        //             15'd406: toneR = `g;     15'd407: toneR = `g;
        //             15'd408: toneR = `g;     15'd409: toneR = `g;
        //             15'd410: toneR = `g;     15'd411: toneR = `g;
        //             15'd412: toneR = `g;     15'd413: toneR = `g;
        //             15'd414: toneR = `g;     15'd415: toneR = `g;
        //             15'd416: toneR = `hc;     15'd417: toneR = `hc;
        //             15'd418: toneR = `hc;     15'd419: toneR = `hc;
        //             15'd420: toneR = `hc;     15'd421: toneR = `hc;
        //             15'd422: toneR = `hc;     15'd423: toneR = `hc;
        //             15'd424: toneR = `hc;     15'd425: toneR = `hc;
        //             15'd426: toneR = `hc;     15'd427: toneR = `hc;
        //             15'd428: toneR = `hc;     15'd429: toneR = `hc;
        //             15'd430: toneR = `hc;     15'd431: toneR = `hc;
        //             15'd432: toneR = `hc;     15'd433: toneR = `hc;
        //             15'd434: toneR = `hc;     15'd435: toneR = `hc;
        //             15'd436: toneR = `hc;     15'd437: toneR = `hc;
        //             15'd438: toneR = `hc;     15'd439: toneR = `hc;
        //             15'd440: toneR = `hc;     15'd441: toneR = `hc;
        //             15'd442: toneR = `hc;     15'd443: toneR = `hc;
        //             15'd444: toneR = `hc;     15'd445: toneR = `hc;
        //             15'd446: toneR = `sil;     15'd447: toneR = `sil;
        //             15'd448: toneR = `hc;     15'd449: toneR = `hc;
        //             15'd450: toneR = `hc;     15'd451: toneR = `hc;
        //             15'd452: toneR = `hc;     15'd453: toneR = `hc;
        //             15'd454: toneR = `hc;     15'd455: toneR = `hc;
        //             15'd456: toneR = `hc;     15'd457: toneR = `hc;
        //             15'd458: toneR = `hc;     15'd459: toneR = `hc;
        //             15'd460: toneR = `hc;     15'd461: toneR = `hc;
        //             15'd462: toneR = `hc;     15'd463: toneR = `hc;
        //             15'd464: toneR = `g;     15'd465: toneR = `g;
        //             15'd466: toneR = `g;     15'd467: toneR = `g;
        //             15'd468: toneR = `g;     15'd469: toneR = `g;
        //             15'd470: toneR = `g;     15'd471: toneR = `g;
        //             15'd472: toneR = `g;     15'd473: toneR = `g;
        //             15'd474: toneR = `g;     15'd475: toneR = `g;
        //             15'd476: toneR = `g;     15'd477: toneR = `g;
        //             15'd478: toneR = `g;     15'd479: toneR = `g;
        //             15'd480: toneR = `hc;     15'd481: toneR = `hc;
        //             15'd482: toneR = `hc;     15'd483: toneR = `hc;
        //             15'd484: toneR = `hc;     15'd485: toneR = `hc;
        //             15'd486: toneR = `hc;     15'd487: toneR = `hc;
        //             15'd488: toneR = `hc;     15'd489: toneR = `hc;
        //             15'd490: toneR = `hc;     15'd491: toneR = `hc;
        //             15'd492: toneR = `hc;     15'd493: toneR = `hc;
        //             15'd494: toneR = `hc;     15'd495: toneR = `hc;
        //             15'd496: toneR = `hc;     15'd497: toneR = `hc;
        //             15'd498: toneR = `hc;     15'd499: toneR = `hc;
        //             15'd500: toneR = `hc;     15'd501: toneR = `hc;
        //             15'd502: toneR = `hc;     15'd503: toneR = `hc;
        //             15'd504: toneR = `hc;     15'd505: toneR = `hc;
        //             15'd506: toneR = `hc;     15'd507: toneR = `hc;
        //             15'd508: toneR = `hc;     15'd509: toneR = `hc;
        //             15'd510: toneR = `hc;     15'd511: toneR = `hc;
        //         default: toneR = `sil;
        //     endcase
         end else begin
             toneR = `sil;
         end
    end

    always @(*) begin
        if(en == 1) begin
            if (_music) begin
                case(ibeatNum)
                    // 15'd0: toneL = `hd;     15'd1: toneL = `hd;
                    // 15'd2: toneL = `hd;     15'd3: toneL = `hd;
                    // 15'd4: toneL = `hd;     15'd5: toneL = `hd;
                    // 15'd6: toneL = `hd;     15'd7: toneL = `hd;
                    // 15'd8: toneL = `hd;     15'd9: toneL = `hd;
                    // 15'd10: toneL = `hd;     15'd11: toneL = `hd;
                    // 15'd12: toneL = `hd;     15'd13: toneL = `hd;
                    // 15'd14: toneL = `hd;     15'd15: toneL = `hd;
                    // 15'd16: toneL = `hd;     15'd17: toneL = `hd;
                    // 15'd18: toneL = `hd;     15'd19: toneL = `hd;
                    // 15'd20: toneL = `hd;     15'd21: toneL = `hd;
                    // 15'd22: toneL = `hd;     15'd23: toneL = `hd;
                    // 15'd24: toneL = `hd;     15'd25: toneL = `hd;
                    // 15'd26: toneL = `hd;     15'd27: toneL = `hd;
                    // 15'd28: toneL = `hd;     15'd29: toneL = `hd;
                    // 15'd30: toneL = `hd;     15'd31: toneL = `hd;
                    // 15'd32: toneL = `a;     15'd33: toneL = `a;
                    // 15'd34: toneL = `a;     15'd35: toneL = `a;
                    // 15'd36: toneL = `a;     15'd37: toneL = `a;
                    // 15'd38: toneL = `a;     15'd39: toneL = `a;
                    // 15'd40: toneL = `a;     15'd41: toneL = `a;
                    // 15'd42: toneL = `a;     15'd43: toneL = `a;
                    // 15'd44: toneL = `a;     15'd45: toneL = `a;
                    // 15'd46: toneL = `a;     15'd47: toneL = `a;
                    // 15'd48: toneL = `a;     15'd49: toneL = `a;
                    // 15'd50: toneL = `a;     15'd51: toneL = `a;
                    // 15'd52: toneL = `a;     15'd53: toneL = `a;
                    // 15'd54: toneL = `a;     15'd55: toneL = `a;
                    // 15'd56: toneL = `a;     15'd57: toneL = `a;
                    // 15'd58: toneL = `a;     15'd59: toneL = `a;
                    // 15'd60: toneL = `a;     15'd61: toneL = `a;
                    // 15'd62: toneL = `a;     15'd63: toneL = `a;
                    // 15'd64: toneL = `b;     15'd65: toneL = `b;
                    // 15'd66: toneL = `b;     15'd67: toneL = `b;
                    // 15'd68: toneL = `b;     15'd69: toneL = `b;
                    // 15'd70: toneL = `b;     15'd71: toneL = `b;
                    // 15'd72: toneL = `b;     15'd73: toneL = `b;
                    // 15'd74: toneL = `b;     15'd75: toneL = `b;
                    // 15'd76: toneL = `b;     15'd77: toneL = `b;
                    // 15'd78: toneL = `b;     15'd79: toneL = `b;
                    // 15'd80: toneL = `b;     15'd81: toneL = `b;
                    // 15'd82: toneL = `b;     15'd83: toneL = `b;
                    // 15'd84: toneL = `b;     15'd85: toneL = `b;
                    // 15'd86: toneL = `b;     15'd87: toneL = `b;
                    // 15'd88: toneL = `b;     15'd89: toneL = `b;
                    // 15'd90: toneL = `b;     15'd91: toneL = `b;
                    // 15'd92: toneL = `b;     15'd93: toneL = `b;
                    // 15'd94: toneL = `b;     15'd95: toneL = `b;
                    // 15'd96: toneL = `rf;     15'd97: toneL = `rf;
                    // 15'd98: toneL = `rf;     15'd99: toneL = `rf;
                    // 15'd100: toneL = `rf;     15'd101: toneL = `rf;
                    // 15'd102: toneL = `rf;     15'd103: toneL = `rf;
                    // 15'd104: toneL = `rf;     15'd105: toneL = `rf;
                    // 15'd106: toneL = `rf;     15'd107: toneL = `rf;
                    // 15'd108: toneL = `rf;     15'd109: toneL = `rf;
                    // 15'd110: toneL = `rf;     15'd111: toneL = `rf;
                    // 15'd112: toneL = `rf;     15'd113: toneL = `rf;
                    // 15'd114: toneL = `rf;     15'd115: toneL = `rf;
                    // 15'd116: toneL = `rf;     15'd117: toneL = `rf;
                    // 15'd118: toneL = `rf;     15'd119: toneL = `rf;
                    // 15'd120: toneL = `rf;     15'd121: toneL = `rf;
                    // 15'd122: toneL = `rf;     15'd123: toneL = `rf;
                    // 15'd124: toneL = `rf;     15'd125: toneL = `rf;
                    // 15'd126: toneL = `rf;     15'd127: toneL = `rf;
                    // 15'd128: toneL = `g;     15'd129: toneL = `g;
                    // 15'd130: toneL = `g;     15'd131: toneL = `g;
                    // 15'd132: toneL = `g;     15'd133: toneL = `g;
                    // 15'd134: toneL = `g;     15'd135: toneL = `g;
                    // 15'd136: toneL = `g;     15'd137: toneL = `g;
                    // 15'd138: toneL = `g;     15'd139: toneL = `g;
                    // 15'd140: toneL = `g;     15'd141: toneL = `g;
                    // 15'd142: toneL = `g;     15'd143: toneL = `g;
                    // 15'd144: toneL = `g;     15'd145: toneL = `g;
                    // 15'd146: toneL = `g;     15'd147: toneL = `g;
                    // 15'd148: toneL = `g;     15'd149: toneL = `g;
                    // 15'd150: toneL = `g;     15'd151: toneL = `g;
                    // 15'd152: toneL = `g;     15'd153: toneL = `g;
                    // 15'd154: toneL = `g;     15'd155: toneL = `g;
                    // 15'd156: toneL = `g;     15'd157: toneL = `g;
                    // 15'd158: toneL = `g;     15'd159: toneL = `g;
                    // 15'd160: toneL = `d;     15'd161: toneL = `d;
                    // 15'd162: toneL = `d;     15'd163: toneL = `d;
                    // 15'd164: toneL = `d;     15'd165: toneL = `d;
                    // 15'd166: toneL = `d;     15'd167: toneL = `d;
                    // 15'd168: toneL = `d;     15'd169: toneL = `d;
                    // 15'd170: toneL = `d;     15'd171: toneL = `d;
                    // 15'd172: toneL = `d;     15'd173: toneL = `d;
                    // 15'd174: toneL = `d;     15'd175: toneL = `d;
                    // 15'd176: toneL = `d;     15'd177: toneL = `d;
                    // 15'd178: toneL = `d;     15'd179: toneL = `d;
                    // 15'd180: toneL = `d;     15'd181: toneL = `d;
                    // 15'd182: toneL = `d;     15'd183: toneL = `d;
                    // 15'd184: toneL = `d;     15'd185: toneL = `d;
                    // 15'd186: toneL = `d;     15'd187: toneL = `d;
                    // 15'd188: toneL = `d;     15'd189: toneL = `d;
                    // 15'd190: toneL = `d;     15'd191: toneL = `d;
                    // 15'd192: toneL = `g;     15'd193: toneL = `g;
                    // 15'd194: toneL = `g;     15'd195: toneL = `g;
                    // 15'd196: toneL = `g;     15'd197: toneL = `g;
                    // 15'd198: toneL = `g;     15'd199: toneL = `g;
                    // 15'd200: toneL = `g;     15'd201: toneL = `g;
                    // 15'd202: toneL = `g;     15'd203: toneL = `g;
                    // 15'd204: toneL = `g;     15'd205: toneL = `g;
                    // 15'd206: toneL = `g;     15'd207: toneL = `g;
                    // 15'd208: toneL = `g;     15'd209: toneL = `g;
                    // 15'd210: toneL = `g;     15'd211: toneL = `g;
                    // 15'd212: toneL = `g;     15'd213: toneL = `g;
                    // 15'd214: toneL = `g;     15'd215: toneL = `g;
                    // 15'd216: toneL = `g;     15'd217: toneL = `g;
                    // 15'd218: toneL = `g;     15'd219: toneL = `g;
                    // 15'd220: toneL = `g;     15'd221: toneL = `g;
                    // 15'd222: toneL = `g;     15'd223: toneL = `g;
                    // 15'd224: toneL = `a;     15'd225: toneL = `a;
                    // 15'd226: toneL = `a;     15'd227: toneL = `a;
                    // 15'd228: toneL = `a;     15'd229: toneL = `a;
                    // 15'd230: toneL = `a;     15'd231: toneL = `a;
                    // 15'd232: toneL = `a;     15'd233: toneL = `a;
                    // 15'd234: toneL = `a;     15'd235: toneL = `a;
                    // 15'd236: toneL = `a;     15'd237: toneL = `a;
                    // 15'd238: toneL = `a;     15'd239: toneL = `a;
                    // 15'd240: toneL = `a;     15'd241: toneL = `a;
                    // 15'd242: toneL = `a;     15'd243: toneL = `a;
                    // 15'd244: toneL = `a;     15'd245: toneL = `a;
                    // 15'd246: toneL = `a;     15'd247: toneL = `a;
                    // 15'd248: toneL = `a;     15'd249: toneL = `a;
                    // 15'd250: toneL = `a;     15'd251: toneL = `a;
                    // 15'd252: toneL = `a;     15'd253: toneL = `a;
                    // 15'd254: toneL = `a;     15'd255: toneL = `a;
                    // 15'd256: toneL = `ha;     15'd257: toneL = `ha;
                    // 15'd258: toneL = `ha;     15'd259: toneL = `ha;
                    // 15'd260: toneL = `ha;     15'd261: toneL = `ha;
                    // 15'd262: toneL = `ha;     15'd263: toneL = `ha;
                    // 15'd264: toneL = `rhf;     15'd265: toneL = `rhf;
                    // 15'd266: toneL = `rhf;     15'd267: toneL = `rhf;
                    // 15'd268: toneL = `hg;     15'd269: toneL = `hg;
                    // 15'd270: toneL = `hg;     15'd271: toneL = `hg;
                    // 15'd272: toneL = `ha;     15'd273: toneL = `ha;
                    // 15'd274: toneL = `ha;     15'd275: toneL = `ha;
                    // 15'd276: toneL = `ha;     15'd277: toneL = `ha;
                    // 15'd278: toneL = `ha;     15'd279: toneL = `ha;
                    // 15'd280: toneL = `rhf;     15'd281: toneL = `rhf;
                    // 15'd282: toneL = `rhf;     15'd283: toneL = `rhf;
                    // 15'd284: toneL = `hg;     15'd285: toneL = `hg;
                    // 15'd286: toneL = `hg;     15'd287: toneL = `hg;
                    // 15'd288: toneL = `ha;     15'd289: toneL = `ha;
                    // 15'd290: toneL = `ha;     15'd291: toneL = `ha;
                    // 15'd292: toneL = `a;     15'd293: toneL = `a;
                    // 15'd294: toneL = `a;     15'd295: toneL = `a;
                    // 15'd296: toneL = `b;     15'd297: toneL = `b;
                    // 15'd298: toneL = `b;     15'd299: toneL = `b;
                    // 15'd300: toneL = `rhc;     15'd301: toneL = `rhc;
                    // 15'd302: toneL = `rhc;     15'd303: toneL = `rhc;
                    // 15'd304: toneL = `hd;     15'd305: toneL = `hd;
                    // 15'd306: toneL = `hd;     15'd307: toneL = `hd;
                    // 15'd308: toneL = `he;     15'd309: toneL = `he;
                    // 15'd310: toneL = `he;     15'd311: toneL = `he;
                    // 15'd312: toneL = `rhf;     15'd313: toneL = `rhf;
                    // 15'd314: toneL = `rhf;     15'd315: toneL = `rhf;
                    // 15'd316: toneL = `hg;     15'd317: toneL = `hg;
                    // 15'd318: toneL = `hg;     15'd319: toneL = `hg;
//                     15'd0: toneL = `sil;     15'd1: toneL = `sil;
// 15'd2: toneL = `sil;     15'd3: toneL = `sil;
// 15'd4: toneL = `sil;     15'd5: toneL = `sil;
// 15'd6: toneL = `sil;     15'd7: toneL = `sil;
// 15'd8: toneL = `a;     15'd9: toneL = `a;
// 15'd10: toneL = `a;     15'd11: toneL = `a;
// 15'd12: toneL = `a;     15'd13: toneL = `a;
// 15'd14: toneL = `a;     15'd15: toneL = `a;
// 15'd16: toneL = `he;     15'd17: toneL = `he;
// 15'd18: toneL = `he;     15'd19: toneL = `he;
// 15'd20: toneL = `he;     15'd21: toneL = `he;
// 15'd22: toneL = `he;     15'd23: toneL = `he;
// 15'd24: toneL = `ha;     15'd25: toneL = `ha;
// 15'd26: toneL = `ha;     15'd27: toneL = `ha;
// 15'd28: toneL = `ha;     15'd29: toneL = `ha;
// 15'd30: toneL = `ha;     15'd31: toneL = `ha;
// 15'd32: toneL = `d;     15'd33: toneL = `d;
// 15'd34: toneL = `d;     15'd35: toneL = `d;
// 15'd36: toneL = `d;     15'd37: toneL = `d;
// 15'd38: toneL = `d;     15'd39: toneL = `d;
// 15'd40: toneL = `a;     15'd41: toneL = `a;
// 15'd42: toneL = `a;     15'd43: toneL = `a;
// 15'd44: toneL = `a;     15'd45: toneL = `a;
// 15'd46: toneL = `a;     15'd47: toneL = `a;
// 15'd48: toneL = `hd;     15'd49: toneL = `hd;
// 15'd50: toneL = `hd;     15'd51: toneL = `hd;
// 15'd52: toneL = `hd;     15'd53: toneL = `hd;
// 15'd54: toneL = `hd;     15'd55: toneL = `hd;
// 15'd56: toneL = `e;     15'd57: toneL = `e;
// 15'd58: toneL = `e;     15'd59: toneL = `e;
// 15'd60: toneL = `e;     15'd61: toneL = `e;
// 15'd62: toneL = `e;     15'd63: toneL = `e;
// 15'd64: toneL = `b;     15'd65: toneL = `b;
// 15'd66: toneL = `b;     15'd67: toneL = `b;
// 15'd68: toneL = `b;     15'd69: toneL = `b;
// 15'd70: toneL = `b;     15'd71: toneL = `b;
// 15'd72: toneL = `he;     15'd73: toneL = `he;
// 15'd74: toneL = `he;     15'd75: toneL = `he;
// 15'd76: toneL = `he;     15'd77: toneL = `he;
// 15'd78: toneL = `he;     15'd79: toneL = `he;
// 15'd80: toneL = `f;     15'd81: toneL = `f;
// 15'd82: toneL = `f;     15'd83: toneL = `f;
// 15'd84: toneL = `f;     15'd85: toneL = `f;
// 15'd86: toneL = `f;     15'd87: toneL = `f;
// 15'd88: toneL = `hc;     15'd89: toneL = `hc;
// 15'd90: toneL = `hc;     15'd91: toneL = `hc;
// 15'd92: toneL = `hc;     15'd93: toneL = `hc;
// 15'd94: toneL = `hc;     15'd95: toneL = `hc;
// 15'd96: toneL = `hf;     15'd97: toneL = `hf;
// 15'd98: toneL = `hf;     15'd99: toneL = `hf;
// 15'd100: toneL = `hf;     15'd101: toneL = `hf;
// 15'd102: toneL = `hf;     15'd103: toneL = `hf;
// 15'd104: toneL = `a;     15'd105: toneL = `a;
// 15'd106: toneL = `a;     15'd107: toneL = `a;
// 15'd108: toneL = `a;     15'd109: toneL = `a;
// 15'd110: toneL = `a;     15'd111: toneL = `a;
// 15'd112: toneL = `he;     15'd113: toneL = `he;
// 15'd114: toneL = `he;     15'd115: toneL = `he;
// 15'd116: toneL = `he;     15'd117: toneL = `he;
// 15'd118: toneL = `he;     15'd119: toneL = `he;
// 15'd120: toneL = `ha;     15'd121: toneL = `ha;
// 15'd122: toneL = `ha;     15'd123: toneL = `ha;
// 15'd124: toneL = `ha;     15'd125: toneL = `ha;
// 15'd126: toneL = `ha;     15'd127: toneL = `ha;
// 15'd128: toneL = `d;     15'd129: toneL = `d;
// 15'd130: toneL = `d;     15'd131: toneL = `d;
// 15'd132: toneL = `d;     15'd133: toneL = `d;
// 15'd134: toneL = `d;     15'd135: toneL = `d;
// 15'd136: toneL = `a;     15'd137: toneL = `a;
// 15'd138: toneL = `a;     15'd139: toneL = `a;
// 15'd140: toneL = `a;     15'd141: toneL = `a;
// 15'd142: toneL = `a;     15'd143: toneL = `a;
// 15'd144: toneL = `hd;     15'd145: toneL = `hd;
// 15'd146: toneL = `hd;     15'd147: toneL = `hd;
// 15'd148: toneL = `hd;     15'd149: toneL = `hd;
// 15'd150: toneL = `hd;     15'd151: toneL = `hd;
// 15'd152: toneL = `e;     15'd153: toneL = `e;
// 15'd154: toneL = `e;     15'd155: toneL = `e;
// 15'd156: toneL = `e;     15'd157: toneL = `e;
// 15'd158: toneL = `e;     15'd159: toneL = `e;
// 15'd160: toneL = `b;     15'd161: toneL = `b;
// 15'd162: toneL = `b;     15'd163: toneL = `b;
// 15'd164: toneL = `b;     15'd165: toneL = `b;
// 15'd166: toneL = `b;     15'd167: toneL = `b;
// 15'd168: toneL = `he;     15'd169: toneL = `he;
// 15'd170: toneL = `he;     15'd171: toneL = `he;
// 15'd172: toneL = `he;     15'd173: toneL = `he;
// 15'd174: toneL = `he;     15'd175: toneL = `he;
// 15'd176: toneL = `a;     15'd177: toneL = `a;
// 15'd178: toneL = `a;     15'd179: toneL = `a;
// 15'd180: toneL = `a;     15'd181: toneL = `a;
// 15'd182: toneL = `a;     15'd183: toneL = `a;
// 15'd184: toneL = `he;     15'd185: toneL = `he;
// 15'd186: toneL = `he;     15'd187: toneL = `he;
// 15'd188: toneL = `he;     15'd189: toneL = `he;
// 15'd190: toneL = `he;     15'd191: toneL = `he;
// 15'd192: toneL = `ha;     15'd193: toneL = `ha;
// 15'd194: toneL = `ha;     15'd195: toneL = `ha;
// 15'd196: toneL = `ha;     15'd197: toneL = `ha;
// 15'd198: toneL = `ha;     15'd199: toneL = `ha;
// 15'd200: toneL = `a;     15'd201: toneL = `a;
// 15'd202: toneL = `a;     15'd203: toneL = `a;
// 15'd204: toneL = `a;     15'd205: toneL = `a;
// 15'd206: toneL = `a;     15'd207: toneL = `a;
// 15'd208: toneL = `he;     15'd209: toneL = `he;
// 15'd210: toneL = `he;     15'd211: toneL = `he;
// 15'd212: toneL = `he;     15'd213: toneL = `he;
// 15'd214: toneL = `he;     15'd215: toneL = `he;
// 15'd216: toneL = `ha;     15'd217: toneL = `ha;
// 15'd218: toneL = `ha;     15'd219: toneL = `ha;
// 15'd220: toneL = `ha;     15'd221: toneL = `ha;
// 15'd222: toneL = `ha;     15'd223: toneL = `ha;
// 15'd224: toneL = `hd;     15'd225: toneL = `hd;
// 15'd226: toneL = `hd;     15'd227: toneL = `hd;
// 15'd228: toneL = `hd;     15'd229: toneL = `hd;
// 15'd230: toneL = `hd;     15'd231: toneL = `hd;
// 15'd232: toneL = `hf;     15'd233: toneL = `hf;
// 15'd234: toneL = `hf;     15'd235: toneL = `hf;
// 15'd236: toneL = `hf;     15'd237: toneL = `hf;
// 15'd238: toneL = `hf;     15'd239: toneL = `hf;
// 15'd240: toneL = `ha;     15'd241: toneL = `ha;
// 15'd242: toneL = `ha;     15'd243: toneL = `ha;
// 15'd244: toneL = `ha;     15'd245: toneL = `ha;
// 15'd246: toneL = `ha;     15'd247: toneL = `ha;
// 15'd248: toneL = `e;     15'd249: toneL = `e;
// 15'd250: toneL = `e;     15'd251: toneL = `e;
// 15'd252: toneL = `e;     15'd253: toneL = `e;
// 15'd254: toneL = `e;     15'd255: toneL = `e;
// 15'd256: toneL = `b;     15'd257: toneL = `b;
// 15'd258: toneL = `b;     15'd259: toneL = `b;
// 15'd260: toneL = `b;     15'd261: toneL = `b;
// 15'd262: toneL = `b;     15'd263: toneL = `b;
// 15'd264: toneL = `he;     15'd265: toneL = `he;
// 15'd266: toneL = `he;     15'd267: toneL = `he;
// 15'd268: toneL = `he;     15'd269: toneL = `he;
// 15'd270: toneL = `he;     15'd271: toneL = `he;
// 15'd272: toneL = `f;     15'd273: toneL = `f;
// 15'd274: toneL = `f;     15'd275: toneL = `f;
// 15'd276: toneL = `f;     15'd277: toneL = `f;
// 15'd278: toneL = `f;     15'd279: toneL = `f;
// 15'd280: toneL = `hc;     15'd281: toneL = `hc;
// 15'd282: toneL = `hc;     15'd283: toneL = `hc;
// 15'd284: toneL = `hc;     15'd285: toneL = `hc;
// 15'd286: toneL = `hc;     15'd287: toneL = `hc;
// 15'd288: toneL = `hf;     15'd289: toneL = `hf;
// 15'd290: toneL = `hf;     15'd291: toneL = `hf;
// 15'd292: toneL = `hf;     15'd293: toneL = `hf;
// 15'd294: toneL = `hf;     15'd295: toneL = `hf;
// 15'd296: toneL = `a;     15'd297: toneL = `a;
// 15'd298: toneL = `a;     15'd299: toneL = `a;
// 15'd300: toneL = `a;     15'd301: toneL = `a;
// 15'd302: toneL = `a;     15'd303: toneL = `a;
// 15'd304: toneL = `he;     15'd305: toneL = `he;
// 15'd306: toneL = `he;     15'd307: toneL = `he;
// 15'd308: toneL = `he;     15'd309: toneL = `he;
// 15'd310: toneL = `he;     15'd311: toneL = `he;
// 15'd312: toneL = `ha;     15'd313: toneL = `ha;
// 15'd314: toneL = `ha;     15'd315: toneL = `ha;
// 15'd316: toneL = `ha;     15'd317: toneL = `ha;
// 15'd318: toneL = `ha;     15'd319: toneL = `ha;
// 15'd320: toneL = `d;     15'd321: toneL = `d;
// 15'd322: toneL = `d;     15'd323: toneL = `d;
// 15'd324: toneL = `d;     15'd325: toneL = `d;
// 15'd326: toneL = `d;     15'd327: toneL = `d;
// 15'd328: toneL = `a;     15'd329: toneL = `a;
// 15'd330: toneL = `a;     15'd331: toneL = `a;
// 15'd332: toneL = `a;     15'd333: toneL = `a;
// 15'd334: toneL = `a;     15'd335: toneL = `a;
// 15'd336: toneL = `hd;     15'd337: toneL = `hd;
// 15'd338: toneL = `hd;     15'd339: toneL = `hd;
// 15'd340: toneL = `hd;     15'd341: toneL = `hd;
// 15'd342: toneL = `hd;     15'd343: toneL = `hd;
// 15'd344: toneL = `e;     15'd345: toneL = `e;
// 15'd346: toneL = `e;     15'd347: toneL = `e;
// 15'd348: toneL = `e;     15'd349: toneL = `e;
// 15'd350: toneL = `e;     15'd351: toneL = `e;
// 15'd352: toneL = `b;     15'd353: toneL = `b;
// 15'd354: toneL = `b;     15'd355: toneL = `b;
// 15'd356: toneL = `b;     15'd357: toneL = `b;
// 15'd358: toneL = `b;     15'd359: toneL = `b;
// 15'd360: toneL = `he;     15'd361: toneL = `he;
// 15'd362: toneL = `he;     15'd363: toneL = `he;
// 15'd364: toneL = `he;     15'd365: toneL = `he;
// 15'd366: toneL = `he;     15'd367: toneL = `he;
// 15'd368: toneL = `a;     15'd369: toneL = `a;
// 15'd370: toneL = `a;     15'd371: toneL = `a;
// 15'd372: toneL = `a;     15'd373: toneL = `a;
// 15'd374: toneL = `a;     15'd375: toneL = `a;
// 15'd376: toneL = `he;     15'd377: toneL = `he;
// 15'd378: toneL = `he;     15'd379: toneL = `he;
// 15'd380: toneL = `he;     15'd381: toneL = `he;
// 15'd382: toneL = `he;     15'd383: toneL = `he;
// 15'd384: toneL = `ha;     15'd385: toneL = `ha;
// 15'd386: toneL = `ha;     15'd387: toneL = `ha;
// 15'd388: toneL = `ha;     15'd389: toneL = `ha;
// 15'd390: toneL = `ha;     15'd391: toneL = `ha;
// 15'd392: toneL = `f;     15'd393: toneL = `f;
// 15'd394: toneL = `f;     15'd395: toneL = `f;
// 15'd396: toneL = `f;     15'd397: toneL = `f;
// 15'd398: toneL = `f;     15'd399: toneL = `f;
// 15'd400: toneL = `hc;     15'd401: toneL = `hc;
// 15'd402: toneL = `hc;     15'd403: toneL = `hc;
// 15'd404: toneL = `hc;     15'd405: toneL = `hc;
// 15'd406: toneL = `hc;     15'd407: toneL = `hc;
// 15'd408: toneL = `hf;     15'd409: toneL = `hf;
// 15'd410: toneL = `hf;     15'd411: toneL = `hf;
// 15'd412: toneL = `hf;     15'd413: toneL = `hf;
// 15'd414: toneL = `hf;     15'd415: toneL = `hf;
// 15'd416: toneL = `e;     15'd417: toneL = `e;
// 15'd418: toneL = `e;     15'd419: toneL = `e;
// 15'd420: toneL = `e;     15'd421: toneL = `e;
// 15'd422: toneL = `e;     15'd423: toneL = `e;
// 15'd424: toneL = `b;     15'd425: toneL = `b;
// 15'd426: toneL = `b;     15'd427: toneL = `b;
// 15'd428: toneL = `b;     15'd429: toneL = `b;
// 15'd430: toneL = `b;     15'd431: toneL = `b;
// 15'd432: toneL = `he;     15'd433: toneL = `he;
// 15'd434: toneL = `he;     15'd435: toneL = `he;
// 15'd436: toneL = `he;     15'd437: toneL = `he;
// 15'd438: toneL = `he;     15'd439: toneL = `he;
// 15'd440: toneL = `a;     15'd441: toneL = `a;
// 15'd442: toneL = `a;     15'd443: toneL = `a;
// 15'd444: toneL = `a;     15'd445: toneL = `a;
// 15'd446: toneL = `a;     15'd447: toneL = `a;
// 15'd448: toneL = `he;     15'd449: toneL = `he;
// 15'd450: toneL = `he;     15'd451: toneL = `he;
// 15'd452: toneL = `he;     15'd453: toneL = `he;
// 15'd454: toneL = `he;     15'd455: toneL = `he;
// 15'd456: toneL = `ha;     15'd457: toneL = `ha;
// 15'd458: toneL = `ha;     15'd459: toneL = `ha;
// 15'd460: toneL = `ha;     15'd461: toneL = `ha;
// 15'd462: toneL = `ha;     15'd463: toneL = `ha;
// 15'd464: toneL = `sil;     15'd465: toneL = `ha;
// 15'd466: toneL = `ha;     15'd467: toneL = `ha;
// 15'd468: toneL = `ha;     15'd469: toneL = `ha;
// 15'd470: toneL = `ha;     15'd471: toneL = `ha;
// 15'd472: toneL = `ha;     15'd473: toneL = `ha;
// 15'd474: toneL = `ha;     15'd475: toneL = `ha;
// 15'd476: toneL = `ha;     15'd477: toneL = `ha;
// 15'd478: toneL = `ha;     15'd479: toneL = `ha;
// 15'd480: toneL = `he;     15'd481: toneL = `he;
// 15'd482: toneL = `he;     15'd483: toneL = `he;
// 15'd484: toneL = `he;     15'd485: toneL = `he;
// 15'd486: toneL = `he;     15'd487: toneL = `he;
// 15'd488: toneL = `ha;     15'd489: toneL = `ha;
// 15'd490: toneL = `ha;     15'd491: toneL = `ha;
// 15'd492: toneL = `ha;     15'd493: toneL = `ha;
// 15'd494: toneL = `ha;     15'd495: toneL = `ha;
// 15'd496: toneL = `hc;     15'd497: toneL = `hc;
// 15'd498: toneL = `hc;     15'd499: toneL = `hc;
// 15'd500: toneL = `hc;     15'd501: toneL = `hc;
// 15'd502: toneL = `hc;     15'd503: toneL = `hc;
// 15'd504: toneL = `a;     15'd505: toneL = `a;
// 15'd506: toneL = `a;     15'd507: toneL = `a;
// 15'd508: toneL = `a;     15'd509: toneL = `a;
// 15'd510: toneL = `a;     15'd511: toneL = `a;
// 15'd512: toneL = `he;     15'd513: toneL = `he;
// 15'd514: toneL = `he;     15'd515: toneL = `he;
// 15'd516: toneL = `he;     15'd517: toneL = `he;
// 15'd518: toneL = `he;     15'd519: toneL = `he;
// 15'd520: toneL = `hb;     15'd521: toneL = `hb;
// 15'd522: toneL = `hb;     15'd523: toneL = `hb;
// 15'd524: toneL = `hb;     15'd525: toneL = `hb;
// 15'd526: toneL = `hb;     15'd527: toneL = `hb;
// 15'd528: toneL = `ha;     15'd529: toneL = `ha;
// 15'd530: toneL = `ha;     15'd531: toneL = `ha;
// 15'd532: toneL = `ha;     15'd533: toneL = `ha;
// 15'd534: toneL = `ha;     15'd535: toneL = `ha;
// 15'd536: toneL = `hhc;     15'd537: toneL = `hhc;
// 15'd538: toneL = `hhc;     15'd539: toneL = `hhc;
// 15'd540: toneL = `hhc;     15'd541: toneL = `hhc;
// 15'd542: toneL = `hhc;     15'd543: toneL = `hhc;
// 15'd544: toneL = `ha;     15'd545: toneL = `ha;
// 15'd546: toneL = `ha;     15'd547: toneL = `ha;
// 15'd548: toneL = `ha;     15'd549: toneL = `ha;
// 15'd550: toneL = `ha;     15'd551: toneL = `ha;
// 15'd552: toneL = `hb;     15'd553: toneL = `hb;
// 15'd554: toneL = `hb;     15'd555: toneL = `hb;
// 15'd556: toneL = `hb;     15'd557: toneL = `hb;
// 15'd558: toneL = `hb;     15'd559: toneL = `hb;
// 15'd560: toneL = `ha;     15'd561: toneL = `ha;
// 15'd562: toneL = `ha;     15'd563: toneL = `ha;
// 15'd564: toneL = `ha;     15'd565: toneL = `ha;
// 15'd566: toneL = `ha;     15'd567: toneL = `ha;
// 15'd568: toneL = `a;     15'd569: toneL = `a;
// 15'd570: toneL = `a;     15'd571: toneL = `a;
// 15'd572: toneL = `a;     15'd573: toneL = `a;
// 15'd574: toneL = `a;     15'd575: toneL = `a;
// 15'd576: toneL = `he;     15'd577: toneL = `he;
// 15'd578: toneL = `he;     15'd579: toneL = `he;
// 15'd580: toneL = `he;     15'd581: toneL = `he;
// 15'd582: toneL = `he;     15'd583: toneL = `he;
// 15'd584: toneL = `ha;     15'd585: toneL = `ha;
// 15'd586: toneL = `ha;     15'd587: toneL = `ha;
// 15'd588: toneL = `ha;     15'd589: toneL = `ha;
// 15'd590: toneL = `ha;     15'd591: toneL = `ha;
// 15'd592: toneL = `hd;     15'd593: toneL = `hd;
// 15'd594: toneL = `hd;     15'd595: toneL = `hd;
// 15'd596: toneL = `hd;     15'd597: toneL = `hd;
// 15'd598: toneL = `hd;     15'd599: toneL = `hd;
// 15'd600: toneL = `hf;     15'd601: toneL = `hf;
// 15'd602: toneL = `hf;     15'd603: toneL = `hf;
// 15'd604: toneL = `hf;     15'd605: toneL = `hf;
// 15'd606: toneL = `hf;     15'd607: toneL = `hf;
// 15'd608: toneL = `ha;     15'd609: toneL = `ha;
// 15'd610: toneL = `ha;     15'd611: toneL = `ha;
// 15'd612: toneL = `ha;     15'd613: toneL = `ha;
// 15'd614: toneL = `ha;     15'd615: toneL = `ha;
// 15'd616: toneL = `e;     15'd617: toneL = `e;
// 15'd618: toneL = `e;     15'd619: toneL = `e;
// 15'd620: toneL = `e;     15'd621: toneL = `e;
// 15'd622: toneL = `e;     15'd623: toneL = `e;
// 15'd624: toneL = `b;     15'd625: toneL = `b;
// 15'd626: toneL = `b;     15'd627: toneL = `b;
// 15'd628: toneL = `b;     15'd629: toneL = `b;
// 15'd630: toneL = `b;     15'd631: toneL = `b;
// 15'd632: toneL = `he;     15'd633: toneL = `he;
// 15'd634: toneL = `he;     15'd635: toneL = `he;
// 15'd636: toneL = `he;     15'd637: toneL = `he;
// 15'd638: toneL = `he;     15'd639: toneL = `he;
// 15'd640: toneL = `f;     15'd641: toneL = `f;
// 15'd642: toneL = `f;     15'd643: toneL = `f;
// 15'd644: toneL = `f;     15'd645: toneL = `f;
// 15'd646: toneL = `f;     15'd647: toneL = `f;
// 15'd648: toneL = `hc;     15'd649: toneL = `hc;
// 15'd650: toneL = `hc;     15'd651: toneL = `hc;
// 15'd652: toneL = `hc;     15'd653: toneL = `hc;
// 15'd654: toneL = `hc;     15'd655: toneL = `hc;
// 15'd656: toneL = `hf;     15'd657: toneL = `hf;
// 15'd658: toneL = `hf;     15'd659: toneL = `hf;
// 15'd660: toneL = `hf;     15'd661: toneL = `hf;
// 15'd662: toneL = `hf;     15'd663: toneL = `hf;
// 15'd664: toneL = `a;     15'd665: toneL = `a;
// 15'd666: toneL = `a;     15'd667: toneL = `a;
// 15'd668: toneL = `a;     15'd669: toneL = `a;
// 15'd670: toneL = `a;     15'd671: toneL = `a;
// 15'd672: toneL = `he;     15'd673: toneL = `he;
// 15'd674: toneL = `he;     15'd675: toneL = `he;
// 15'd676: toneL = `he;     15'd677: toneL = `he;
// 15'd678: toneL = `he;     15'd679: toneL = `he;
// 15'd680: toneL = `ha;     15'd681: toneL = `ha;
// 15'd682: toneL = `ha;     15'd683: toneL = `ha;
// 15'd684: toneL = `ha;     15'd685: toneL = `ha;
// 15'd686: toneL = `ha;     15'd687: toneL = `ha;
// 15'd688: toneL = `d;     15'd689: toneL = `d;
// 15'd690: toneL = `d;     15'd691: toneL = `d;
// 15'd692: toneL = `d;     15'd693: toneL = `d;
// 15'd694: toneL = `d;     15'd695: toneL = `d;
// 15'd696: toneL = `a;     15'd697: toneL = `a;
// 15'd698: toneL = `a;     15'd699: toneL = `a;
// 15'd700: toneL = `a;     15'd701: toneL = `a;
// 15'd702: toneL = `a;     15'd703: toneL = `a;
// 15'd704: toneL = `hd;     15'd705: toneL = `hd;
// 15'd706: toneL = `hd;     15'd707: toneL = `hd;
// 15'd708: toneL = `hd;     15'd709: toneL = `hd;
// 15'd710: toneL = `hd;     15'd711: toneL = `hd;
// 15'd712: toneL = `e;     15'd713: toneL = `e;
// 15'd714: toneL = `e;     15'd715: toneL = `e;
// 15'd716: toneL = `e;     15'd717: toneL = `e;
// 15'd718: toneL = `e;     15'd719: toneL = `e;
// 15'd720: toneL = `b;     15'd721: toneL = `b;
// 15'd722: toneL = `b;     15'd723: toneL = `b;
// 15'd724: toneL = `b;     15'd725: toneL = `b;
// 15'd726: toneL = `b;     15'd727: toneL = `b;
// 15'd728: toneL = `he;     15'd729: toneL = `he;
// 15'd730: toneL = `he;     15'd731: toneL = `he;
// 15'd732: toneL = `he;     15'd733: toneL = `he;
// 15'd734: toneL = `he;     15'd735: toneL = `he;
// 15'd736: toneL = `a;     15'd737: toneL = `a;
// 15'd738: toneL = `a;     15'd739: toneL = `a;
// 15'd740: toneL = `a;     15'd741: toneL = `a;
// 15'd742: toneL = `a;     15'd743: toneL = `a;
// 15'd744: toneL = `he;     15'd745: toneL = `he;
// 15'd746: toneL = `he;     15'd747: toneL = `he;
// 15'd748: toneL = `he;     15'd749: toneL = `he;
// 15'd750: toneL = `he;     15'd751: toneL = `he;
// 15'd752: toneL = `ha;     15'd753: toneL = `ha;
// 15'd754: toneL = `ha;     15'd755: toneL = `ha;
// 15'd756: toneL = `ha;     15'd757: toneL = `ha;
// 15'd758: toneL = `ha;     15'd759: toneL = `ha;
// 15'd760: toneL = `f;     15'd761: toneL = `f;
// 15'd762: toneL = `f;     15'd763: toneL = `f;
// 15'd764: toneL = `f;     15'd765: toneL = `f;
// 15'd766: toneL = `f;     15'd767: toneL = `f;
// 15'd768: toneL = `hc;     15'd769: toneL = `hc;
// 15'd770: toneL = `hc;     15'd771: toneL = `hc;
// 15'd772: toneL = `hc;     15'd773: toneL = `hc;
// 15'd774: toneL = `hc;     15'd775: toneL = `hc;
// 15'd776: toneL = `hf;     15'd777: toneL = `hf;
// 15'd778: toneL = `hf;     15'd779: toneL = `hf;
// 15'd780: toneL = `hf;     15'd781: toneL = `hf;
// 15'd782: toneL = `hf;     15'd783: toneL = `hf;
// 15'd784: toneL = `e;     15'd785: toneL = `e;
// 15'd786: toneL = `e;     15'd787: toneL = `e;
// 15'd788: toneL = `e;     15'd789: toneL = `e;
// 15'd790: toneL = `e;     15'd791: toneL = `e;
// 15'd792: toneL = `b;     15'd793: toneL = `b;
// 15'd794: toneL = `b;     15'd795: toneL = `b;
// 15'd796: toneL = `b;     15'd797: toneL = `b;
// 15'd798: toneL = `b;     15'd799: toneL = `b;
// 15'd800: toneL = `he;     15'd801: toneL = `he;
// 15'd802: toneL = `he;     15'd803: toneL = `he;
// 15'd804: toneL = `he;     15'd805: toneL = `he;
// 15'd806: toneL = `he;     15'd807: toneL = `he;
15'd0: toneL = `sil;     15'd1: toneL = `sil;
15'd2: toneL = `sil;     15'd3: toneL = `sil;
15'd4: toneL = `sil;     15'd5: toneL = `sil;
15'd6: toneL = `sil;     15'd7: toneL = `sil;
15'd8: toneL = `a;     15'd9: toneL = `a;
15'd10: toneL = `a;     15'd11: toneL = `a;
15'd12: toneL = `a;     15'd13: toneL = `a;
15'd14: toneL = `a;     15'd15: toneL = `a;
15'd16: toneL = `he;     15'd17: toneL = `he;
15'd18: toneL = `he;     15'd19: toneL = `he;
15'd20: toneL = `he;     15'd21: toneL = `he;
15'd22: toneL = `he;     15'd23: toneL = `he;
15'd24: toneL = `ha;     15'd25: toneL = `ha;
15'd26: toneL = `ha;     15'd27: toneL = `ha;
15'd28: toneL = `ha;     15'd29: toneL = `ha;
15'd30: toneL = `ha;     15'd31: toneL = `ha;
15'd32: toneL = `ha;     15'd33: toneL = `ha;
15'd34: toneL = `ha;     15'd35: toneL = `ha;
15'd36: toneL = `ha;     15'd37: toneL = `ha;
15'd38: toneL = `ha;     15'd39: toneL = `ha;
15'd40: toneL = `d;     15'd41: toneL = `d;
15'd42: toneL = `d;     15'd43: toneL = `d;
15'd44: toneL = `d;     15'd45: toneL = `d;
15'd46: toneL = `d;     15'd47: toneL = `d;
15'd48: toneL = `a;     15'd49: toneL = `a;
15'd50: toneL = `a;     15'd51: toneL = `a;
15'd52: toneL = `a;     15'd53: toneL = `a;
15'd54: toneL = `a;     15'd55: toneL = `a;
15'd56: toneL = `hd;     15'd57: toneL = `hd;
15'd58: toneL = `hd;     15'd59: toneL = `hd;
15'd60: toneL = `hd;     15'd61: toneL = `hd;
15'd62: toneL = `hd;     15'd63: toneL = `hd;
15'd64: toneL = `hd;     15'd65: toneL = `hd;
15'd66: toneL = `hd;     15'd67: toneL = `hd;
15'd68: toneL = `hd;     15'd69: toneL = `hd;
15'd70: toneL = `hd;     15'd71: toneL = `hd;
15'd72: toneL = `e;     15'd73: toneL = `e;
15'd74: toneL = `e;     15'd75: toneL = `e;
15'd76: toneL = `e;     15'd77: toneL = `e;
15'd78: toneL = `e;     15'd79: toneL = `e;
15'd80: toneL = `b;     15'd81: toneL = `b;
15'd82: toneL = `b;     15'd83: toneL = `b;
15'd84: toneL = `b;     15'd85: toneL = `b;
15'd86: toneL = `b;     15'd87: toneL = `b;
15'd88: toneL = `he;     15'd89: toneL = `he;
15'd90: toneL = `he;     15'd91: toneL = `he;
15'd92: toneL = `he;     15'd93: toneL = `he;
15'd94: toneL = `he;     15'd95: toneL = `he;
15'd96: toneL = `he;     15'd97: toneL = `he;
15'd98: toneL = `he;     15'd99: toneL = `he;
15'd100: toneL = `he;     15'd101: toneL = `he;
15'd102: toneL = `he;     15'd103: toneL = `he;
15'd104: toneL = `f;     15'd105: toneL = `f;
15'd106: toneL = `f;     15'd107: toneL = `f;
15'd108: toneL = `f;     15'd109: toneL = `f;
15'd110: toneL = `f;     15'd111: toneL = `f;
15'd112: toneL = `hc;     15'd113: toneL = `hc;
15'd114: toneL = `hc;     15'd115: toneL = `hc;
15'd116: toneL = `hc;     15'd117: toneL = `hc;
15'd118: toneL = `hc;     15'd119: toneL = `hc;
15'd120: toneL = `hf;     15'd121: toneL = `hf;
15'd122: toneL = `hf;     15'd123: toneL = `hf;
15'd124: toneL = `hf;     15'd125: toneL = `hf;
15'd126: toneL = `hf;     15'd127: toneL = `hf;
15'd128: toneL = `hf;     15'd129: toneL = `hf;
15'd130: toneL = `hf;     15'd131: toneL = `hf;
15'd132: toneL = `hf;     15'd133: toneL = `hf;
15'd134: toneL = `hf;     15'd135: toneL = `hf;
15'd136: toneL = `a;     15'd137: toneL = `a;
15'd138: toneL = `a;     15'd139: toneL = `a;
15'd140: toneL = `a;     15'd141: toneL = `a;
15'd142: toneL = `a;     15'd143: toneL = `a;
15'd144: toneL = `hc;     15'd145: toneL = `hc;
15'd146: toneL = `hc;     15'd147: toneL = `hc;
15'd148: toneL = `hc;     15'd149: toneL = `hc;
15'd150: toneL = `hc;     15'd151: toneL = `hc;
15'd152: toneL = `ha;     15'd153: toneL = `ha;
15'd154: toneL = `ha;     15'd155: toneL = `ha;
15'd156: toneL = `ha;     15'd157: toneL = `ha;
15'd158: toneL = `ha;     15'd159: toneL = `ha;
15'd160: toneL = `ha;     15'd161: toneL = `ha;
15'd162: toneL = `ha;     15'd163: toneL = `ha;
15'd164: toneL = `ha;     15'd165: toneL = `ha;
15'd166: toneL = `ha;     15'd167: toneL = `ha;
15'd168: toneL = `d;     15'd169: toneL = `d;
15'd170: toneL = `d;     15'd171: toneL = `d;
15'd172: toneL = `d;     15'd173: toneL = `d;
15'd174: toneL = `d;     15'd175: toneL = `d;
15'd176: toneL = `a;     15'd177: toneL = `a;
15'd178: toneL = `a;     15'd179: toneL = `a;
15'd180: toneL = `a;     15'd181: toneL = `a;
15'd182: toneL = `a;     15'd183: toneL = `a;
15'd184: toneL = `hd;     15'd185: toneL = `hd;
15'd186: toneL = `hd;     15'd187: toneL = `hd;
15'd188: toneL = `hd;     15'd189: toneL = `hd;
15'd190: toneL = `hd;     15'd191: toneL = `hd;
15'd192: toneL = `hd;     15'd193: toneL = `hd;
15'd194: toneL = `hd;     15'd195: toneL = `hd;
15'd196: toneL = `hd;     15'd197: toneL = `hd;
15'd198: toneL = `hd;     15'd199: toneL = `hd;
15'd200: toneL = `e;     15'd201: toneL = `e;
15'd202: toneL = `e;     15'd203: toneL = `e;
15'd204: toneL = `e;     15'd205: toneL = `e;
15'd206: toneL = `e;     15'd207: toneL = `e;
15'd208: toneL = `b;     15'd209: toneL = `b;
15'd210: toneL = `b;     15'd211: toneL = `b;
15'd212: toneL = `b;     15'd213: toneL = `b;
15'd214: toneL = `b;     15'd215: toneL = `b;
15'd216: toneL = `he;     15'd217: toneL = `he;
15'd218: toneL = `he;     15'd219: toneL = `he;
15'd220: toneL = `he;     15'd221: toneL = `he;
15'd222: toneL = `he;     15'd223: toneL = `he;
15'd224: toneL = `he;     15'd225: toneL = `he;
15'd226: toneL = `he;     15'd227: toneL = `he;
15'd228: toneL = `he;     15'd229: toneL = `he;
15'd230: toneL = `he;     15'd231: toneL = `he;
15'd232: toneL = `a;     15'd233: toneL = `a;
15'd234: toneL = `a;     15'd235: toneL = `a;
15'd236: toneL = `a;     15'd237: toneL = `a;
15'd238: toneL = `a;     15'd239: toneL = `a;
15'd240: toneL = `he;     15'd241: toneL = `he;
15'd242: toneL = `he;     15'd243: toneL = `he;
15'd244: toneL = `he;     15'd245: toneL = `he;
15'd246: toneL = `he;     15'd247: toneL = `he;
15'd248: toneL = `ha;     15'd249: toneL = `ha;
15'd250: toneL = `ha;     15'd251: toneL = `ha;
15'd252: toneL = `ha;     15'd253: toneL = `ha;
15'd254: toneL = `ha;     15'd255: toneL = `ha;
15'd256: toneL = `ha;     15'd257: toneL = `ha;
15'd258: toneL = `ha;     15'd259: toneL = `ha;
15'd260: toneL = `ha;     15'd261: toneL = `ha;
15'd262: toneL = `ha;     15'd263: toneL = `ha;
15'd264: toneL = `a;     15'd265: toneL = `a;
15'd266: toneL = `a;     15'd267: toneL = `a;
15'd268: toneL = `a;     15'd269: toneL = `a;
15'd270: toneL = `a;     15'd271: toneL = `a;
15'd272: toneL = `hc;     15'd273: toneL = `hc;
15'd274: toneL = `hc;     15'd275: toneL = `hc;
15'd276: toneL = `hc;     15'd277: toneL = `hc;
15'd278: toneL = `hc;     15'd279: toneL = `hc;
15'd280: toneL = `ha;     15'd281: toneL = `ha;
15'd282: toneL = `ha;     15'd283: toneL = `ha;
15'd284: toneL = `ha;     15'd285: toneL = `ha;
15'd286: toneL = `ha;     15'd287: toneL = `ha;
15'd288: toneL = `ha;     15'd289: toneL = `ha;
15'd290: toneL = `ha;     15'd291: toneL = `ha;
15'd292: toneL = `ha;     15'd293: toneL = `ha;
15'd294: toneL = `ha;     15'd295: toneL = `ha;
15'd296: toneL = `hd;     15'd297: toneL = `hd;
15'd298: toneL = `hd;     15'd299: toneL = `hd;
15'd300: toneL = `hd;     15'd301: toneL = `hd;
15'd302: toneL = `hd;     15'd303: toneL = `hd;
15'd304: toneL = `hf;     15'd305: toneL = `hf;
15'd306: toneL = `hf;     15'd307: toneL = `hf;
15'd308: toneL = `hf;     15'd309: toneL = `hf;
15'd310: toneL = `hf;     15'd311: toneL = `hf;
15'd312: toneL = `ha;     15'd313: toneL = `ha;
15'd314: toneL = `ha;     15'd315: toneL = `ha;
15'd316: toneL = `ha;     15'd317: toneL = `ha;
15'd318: toneL = `ha;     15'd319: toneL = `ha;
15'd320: toneL = `ha;     15'd321: toneL = `ha;
15'd322: toneL = `ha;     15'd323: toneL = `ha;
15'd324: toneL = `ha;     15'd325: toneL = `ha;
15'd326: toneL = `ha;     15'd327: toneL = `ha;
15'd328: toneL = `e;     15'd329: toneL = `e;
15'd330: toneL = `e;     15'd331: toneL = `e;
15'd332: toneL = `e;     15'd333: toneL = `e;
15'd334: toneL = `e;     15'd335: toneL = `e;
15'd336: toneL = `b;     15'd337: toneL = `b;
15'd338: toneL = `b;     15'd339: toneL = `b;
15'd340: toneL = `b;     15'd341: toneL = `b;
15'd342: toneL = `b;     15'd343: toneL = `b;
15'd344: toneL = `he;     15'd345: toneL = `he;
15'd346: toneL = `he;     15'd347: toneL = `he;
15'd348: toneL = `he;     15'd349: toneL = `he;
15'd350: toneL = `he;     15'd351: toneL = `he;
15'd352: toneL = `he;     15'd353: toneL = `he;
15'd354: toneL = `he;     15'd355: toneL = `he;
15'd356: toneL = `he;     15'd357: toneL = `he;
15'd358: toneL = `he;     15'd359: toneL = `he;
15'd360: toneL = `f;     15'd361: toneL = `f;
15'd362: toneL = `f;     15'd363: toneL = `f;
15'd364: toneL = `f;     15'd365: toneL = `f;
15'd366: toneL = `f;     15'd367: toneL = `f;
15'd368: toneL = `hc;     15'd369: toneL = `hc;
15'd370: toneL = `hc;     15'd371: toneL = `hc;
15'd372: toneL = `hc;     15'd373: toneL = `hc;
15'd374: toneL = `hc;     15'd375: toneL = `hc;
15'd376: toneL = `hf;     15'd377: toneL = `hf;
15'd378: toneL = `hf;     15'd379: toneL = `hf;
15'd380: toneL = `hf;     15'd381: toneL = `hf;
15'd382: toneL = `hf;     15'd383: toneL = `hf;
15'd384: toneL = `hf;     15'd385: toneL = `hf;
15'd386: toneL = `hf;     15'd387: toneL = `hf;
15'd388: toneL = `hf;     15'd389: toneL = `hf;
15'd390: toneL = `hf;     15'd391: toneL = `hf;
15'd392: toneL = `a;     15'd393: toneL = `a;
15'd394: toneL = `a;     15'd395: toneL = `a;
15'd396: toneL = `a;     15'd397: toneL = `a;
15'd398: toneL = `a;     15'd399: toneL = `a;
15'd400: toneL = `hc;     15'd401: toneL = `hc;
15'd402: toneL = `hc;     15'd403: toneL = `hc;
15'd404: toneL = `hc;     15'd405: toneL = `hc;
15'd406: toneL = `hc;     15'd407: toneL = `hc;
15'd408: toneL = `ha;     15'd409: toneL = `ha;
15'd410: toneL = `ha;     15'd411: toneL = `ha;
15'd412: toneL = `ha;     15'd413: toneL = `ha;
15'd414: toneL = `ha;     15'd415: toneL = `ha;
15'd416: toneL = `ha;     15'd417: toneL = `ha;
15'd418: toneL = `ha;     15'd419: toneL = `ha;
15'd420: toneL = `ha;     15'd421: toneL = `ha;
15'd422: toneL = `ha;     15'd423: toneL = `ha;
15'd424: toneL = `d;     15'd425: toneL = `d;
15'd426: toneL = `d;     15'd427: toneL = `d;
15'd428: toneL = `d;     15'd429: toneL = `d;
15'd430: toneL = `d;     15'd431: toneL = `d;
15'd432: toneL = `a;     15'd433: toneL = `a;
15'd434: toneL = `a;     15'd435: toneL = `a;
15'd436: toneL = `a;     15'd437: toneL = `a;
15'd438: toneL = `a;     15'd439: toneL = `a;
15'd440: toneL = `hd;     15'd441: toneL = `hd;
15'd442: toneL = `hd;     15'd443: toneL = `hd;
15'd444: toneL = `hd;     15'd445: toneL = `hd;
15'd446: toneL = `hd;     15'd447: toneL = `hd;
15'd448: toneL = `hd;     15'd449: toneL = `hd;
15'd450: toneL = `hd;     15'd451: toneL = `hd;
15'd452: toneL = `hd;     15'd453: toneL = `hd;
15'd454: toneL = `hd;     15'd455: toneL = `hd;
15'd456: toneL = `e;     15'd457: toneL = `e;
15'd458: toneL = `e;     15'd459: toneL = `e;
15'd460: toneL = `e;     15'd461: toneL = `e;
15'd462: toneL = `e;     15'd463: toneL = `e;
15'd464: toneL = `b;     15'd465: toneL = `b;
15'd466: toneL = `b;     15'd467: toneL = `b;
15'd468: toneL = `b;     15'd469: toneL = `b;
15'd470: toneL = `b;     15'd471: toneL = `b;
15'd472: toneL = `he;     15'd473: toneL = `he;
15'd474: toneL = `he;     15'd475: toneL = `he;
15'd476: toneL = `he;     15'd477: toneL = `he;
15'd478: toneL = `he;     15'd479: toneL = `he;
15'd480: toneL = `he;     15'd481: toneL = `he;
15'd482: toneL = `he;     15'd483: toneL = `he;
15'd484: toneL = `he;     15'd485: toneL = `he;
15'd486: toneL = `he;     15'd487: toneL = `he;
15'd488: toneL = `a;     15'd489: toneL = `a;
15'd490: toneL = `a;     15'd491: toneL = `a;
15'd492: toneL = `a;     15'd493: toneL = `a;
15'd494: toneL = `a;     15'd495: toneL = `a;
15'd496: toneL = `he;     15'd497: toneL = `he;
15'd498: toneL = `he;     15'd499: toneL = `he;
15'd500: toneL = `he;     15'd501: toneL = `he;
15'd502: toneL = `he;     15'd503: toneL = `he;
15'd504: toneL = `ha;     15'd505: toneL = `ha;
15'd506: toneL = `ha;     15'd507: toneL = `ha;
15'd508: toneL = `ha;     15'd509: toneL = `ha;
15'd510: toneL = `ha;     15'd511: toneL = `ha;
15'd512: toneL = `ha;     15'd513: toneL = `ha;
15'd514: toneL = `ha;     15'd515: toneL = `ha;
15'd516: toneL = `ha;     15'd517: toneL = `ha;
15'd518: toneL = `ha;     15'd519: toneL = `ha;
15'd520: toneL = `f;     15'd521: toneL = `f;
15'd522: toneL = `f;     15'd523: toneL = `f;
15'd524: toneL = `f;     15'd525: toneL = `f;
15'd526: toneL = `f;     15'd527: toneL = `f;
15'd528: toneL = `hc;     15'd529: toneL = `hc;
15'd530: toneL = `hc;     15'd531: toneL = `hc;
15'd532: toneL = `hc;     15'd533: toneL = `hc;
15'd534: toneL = `hc;     15'd535: toneL = `hc;
15'd536: toneL = `hf;     15'd537: toneL = `hf;
15'd538: toneL = `hf;     15'd539: toneL = `hf;
15'd540: toneL = `hf;     15'd541: toneL = `hf;
15'd542: toneL = `hf;     15'd543: toneL = `hf;
15'd544: toneL = `hf;     15'd545: toneL = `hf;
15'd546: toneL = `hf;     15'd547: toneL = `hf;
15'd548: toneL = `hf;     15'd549: toneL = `hf;
15'd550: toneL = `hf;     15'd551: toneL = `hf;
15'd552: toneL = `e;     15'd553: toneL = `e;
15'd554: toneL = `e;     15'd555: toneL = `e;
15'd556: toneL = `e;     15'd557: toneL = `e;
15'd558: toneL = `e;     15'd559: toneL = `e;
15'd560: toneL = `b;     15'd561: toneL = `b;
15'd562: toneL = `b;     15'd563: toneL = `b;
15'd564: toneL = `b;     15'd565: toneL = `b;
15'd566: toneL = `b;     15'd567: toneL = `b;
15'd568: toneL = `he;     15'd569: toneL = `he;
15'd570: toneL = `he;     15'd571: toneL = `he;
15'd572: toneL = `he;     15'd573: toneL = `he;
15'd574: toneL = `he;     15'd575: toneL = `he;
15'd576: toneL = `he;     15'd577: toneL = `he;
15'd578: toneL = `he;     15'd579: toneL = `he;
15'd580: toneL = `he;     15'd581: toneL = `he;
15'd582: toneL = `he;     15'd583: toneL = `he;
15'd584: toneL = `a;     15'd585: toneL = `a;
15'd586: toneL = `a;     15'd587: toneL = `a;
15'd588: toneL = `a;     15'd589: toneL = `a;
15'd590: toneL = `a;     15'd591: toneL = `a;
15'd592: toneL = `he;     15'd593: toneL = `he;
15'd594: toneL = `he;     15'd595: toneL = `he;
15'd596: toneL = `he;     15'd597: toneL = `he;
15'd598: toneL = `he;     15'd599: toneL = `he;
15'd600: toneL = `ha;     15'd601: toneL = `ha;
15'd602: toneL = `ha;     15'd603: toneL = `ha;
15'd604: toneL = `ha;     15'd605: toneL = `ha;
15'd606: toneL = `ha;     15'd607: toneL = `ha;
15'd608: toneL = `sil;     15'd609: toneL = `ha;
15'd610: toneL = `ha;     15'd611: toneL = `ha;
15'd612: toneL = `ha;     15'd613: toneL = `ha;
15'd614: toneL = `ha;     15'd615: toneL = `ha;
15'd616: toneL = `he;     15'd617: toneL = `he;
15'd618: toneL = `he;     15'd619: toneL = `he;
15'd620: toneL = `he;     15'd621: toneL = `he;
15'd622: toneL = `he;     15'd623: toneL = `he;
15'd624: toneL = `ha;     15'd625: toneL = `ha;
15'd626: toneL = `ha;     15'd627: toneL = `ha;
15'd628: toneL = `ha;     15'd629: toneL = `ha;
15'd630: toneL = `ha;     15'd631: toneL = `ha;
15'd632: toneL = `he;     15'd633: toneL = `he;
15'd634: toneL = `he;     15'd635: toneL = `he;
15'd636: toneL = `he;     15'd637: toneL = `he;
15'd638: toneL = `he;     15'd639: toneL = `he;
15'd640: toneL = `a;     15'd641: toneL = `a;
15'd642: toneL = `a;     15'd643: toneL = `a;
15'd644: toneL = `a;     15'd645: toneL = `a;
15'd646: toneL = `a;     15'd647: toneL = `a;
15'd648: toneL = `he;     15'd649: toneL = `he;
15'd650: toneL = `he;     15'd651: toneL = `he;
15'd652: toneL = `he;     15'd653: toneL = `he;
15'd654: toneL = `he;     15'd655: toneL = `he;
15'd656: toneL = `hb;     15'd657: toneL = `hb;
15'd658: toneL = `hb;     15'd659: toneL = `hb;
15'd660: toneL = `hb;     15'd661: toneL = `hb;
15'd662: toneL = `hb;     15'd663: toneL = `hb;
15'd664: toneL = `ha;     15'd665: toneL = `ha;
15'd666: toneL = `ha;     15'd667: toneL = `ha;
15'd668: toneL = `ha;     15'd669: toneL = `ha;
15'd670: toneL = `ha;     15'd671: toneL = `ha;
15'd672: toneL = `hhc;     15'd673: toneL = `hhc;
15'd674: toneL = `hhc;     15'd675: toneL = `hhc;
15'd676: toneL = `hhc;     15'd677: toneL = `hhc;
15'd678: toneL = `hhc;     15'd679: toneL = `hhc;
15'd680: toneL = `ha;     15'd681: toneL = `ha;
15'd682: toneL = `ha;     15'd683: toneL = `ha;
15'd684: toneL = `ha;     15'd685: toneL = `ha;
15'd686: toneL = `ha;     15'd687: toneL = `ha;
15'd688: toneL = `hb;     15'd689: toneL = `hb;
15'd690: toneL = `hb;     15'd691: toneL = `hb;
15'd692: toneL = `hb;     15'd693: toneL = `hb;
15'd694: toneL = `hb;     15'd695: toneL = `hb;
15'd696: toneL = `ha;     15'd697: toneL = `ha;
15'd698: toneL = `ha;     15'd699: toneL = `ha;
15'd700: toneL = `ha;     15'd701: toneL = `ha;
15'd702: toneL = `ha;     15'd703: toneL = `ha;
15'd704: toneL = `a;     15'd705: toneL = `a;
15'd706: toneL = `a;     15'd707: toneL = `a;
15'd708: toneL = `a;     15'd709: toneL = `a;
15'd710: toneL = `a;     15'd711: toneL = `a;
15'd712: toneL = `he;     15'd713: toneL = `he;
15'd714: toneL = `he;     15'd715: toneL = `he;
15'd716: toneL = `he;     15'd717: toneL = `he;
15'd718: toneL = `he;     15'd719: toneL = `he;
15'd720: toneL = `ha;     15'd721: toneL = `ha;
15'd722: toneL = `ha;     15'd723: toneL = `ha;
15'd724: toneL = `ha;     15'd725: toneL = `ha;
15'd726: toneL = `ha;     15'd727: toneL = `ha;
15'd728: toneL = `ha;     15'd729: toneL = `ha;
15'd730: toneL = `ha;     15'd731: toneL = `ha;
15'd732: toneL = `ha;     15'd733: toneL = `ha;
15'd734: toneL = `ha;     15'd735: toneL = `ha;
15'd736: toneL = `hd;     15'd737: toneL = `hd;
15'd738: toneL = `hd;     15'd739: toneL = `hd;
15'd740: toneL = `hd;     15'd741: toneL = `hd;
15'd742: toneL = `hd;     15'd743: toneL = `hd;
15'd744: toneL = `hf;     15'd745: toneL = `hf;
15'd746: toneL = `hf;     15'd747: toneL = `hf;
15'd748: toneL = `hf;     15'd749: toneL = `hf;
15'd750: toneL = `hf;     15'd751: toneL = `hf;
15'd752: toneL = `ha;     15'd753: toneL = `ha;
15'd754: toneL = `ha;     15'd755: toneL = `ha;
15'd756: toneL = `ha;     15'd757: toneL = `ha;
15'd758: toneL = `ha;     15'd759: toneL = `ha;
15'd760: toneL = `ha;     15'd761: toneL = `ha;
15'd762: toneL = `ha;     15'd763: toneL = `ha;
15'd764: toneL = `ha;     15'd765: toneL = `ha;
15'd766: toneL = `ha;     15'd767: toneL = `ha;
15'd768: toneL = `e;     15'd769: toneL = `e;
15'd770: toneL = `e;     15'd771: toneL = `e;
15'd772: toneL = `e;     15'd773: toneL = `e;
15'd774: toneL = `e;     15'd775: toneL = `e;
15'd776: toneL = `b;     15'd777: toneL = `b;
15'd778: toneL = `b;     15'd779: toneL = `b;
15'd780: toneL = `b;     15'd781: toneL = `b;
15'd782: toneL = `b;     15'd783: toneL = `b;
15'd784: toneL = `he;     15'd785: toneL = `he;
15'd786: toneL = `he;     15'd787: toneL = `he;
15'd788: toneL = `he;     15'd789: toneL = `he;
15'd790: toneL = `he;     15'd791: toneL = `he;
15'd792: toneL = `he;     15'd793: toneL = `he;
15'd794: toneL = `he;     15'd795: toneL = `he;
15'd796: toneL = `he;     15'd797: toneL = `he;
15'd798: toneL = `he;     15'd799: toneL = `he;
15'd800: toneL = `f;     15'd801: toneL = `f;
15'd802: toneL = `f;     15'd803: toneL = `f;
15'd804: toneL = `f;     15'd805: toneL = `f;
15'd806: toneL = `f;     15'd807: toneL = `f;
15'd808: toneL = `hc;     15'd809: toneL = `hc;
15'd810: toneL = `hc;     15'd811: toneL = `hc;
15'd812: toneL = `hc;     15'd813: toneL = `hc;
15'd814: toneL = `hc;     15'd815: toneL = `hc;
15'd816: toneL = `hf;     15'd817: toneL = `hf;
15'd818: toneL = `hf;     15'd819: toneL = `hf;
15'd820: toneL = `hf;     15'd821: toneL = `hf;
15'd822: toneL = `hf;     15'd823: toneL = `hf;
15'd824: toneL = `hf;     15'd825: toneL = `hf;
15'd826: toneL = `hf;     15'd827: toneL = `hf;
15'd828: toneL = `hf;     15'd829: toneL = `hf;
15'd830: toneL = `hf;     15'd831: toneL = `hf;
15'd832: toneL = `a;     15'd833: toneL = `a;
15'd834: toneL = `a;     15'd835: toneL = `a;
15'd836: toneL = `a;     15'd837: toneL = `a;
15'd838: toneL = `a;     15'd839: toneL = `a;
15'd840: toneL = `hc;     15'd841: toneL = `hc;
15'd842: toneL = `hc;     15'd843: toneL = `hc;
15'd844: toneL = `hc;     15'd845: toneL = `hc;
15'd846: toneL = `hc;     15'd847: toneL = `hc;
15'd848: toneL = `ha;     15'd849: toneL = `ha;
15'd850: toneL = `ha;     15'd851: toneL = `ha;
15'd852: toneL = `ha;     15'd853: toneL = `ha;
15'd854: toneL = `ha;     15'd855: toneL = `ha;
15'd856: toneL = `ha;     15'd857: toneL = `ha;
15'd858: toneL = `ha;     15'd859: toneL = `ha;
15'd860: toneL = `ha;     15'd861: toneL = `ha;
15'd862: toneL = `ha;     15'd863: toneL = `ha;
15'd864: toneL = `d;     15'd865: toneL = `d;
15'd866: toneL = `d;     15'd867: toneL = `d;
15'd868: toneL = `d;     15'd869: toneL = `d;
15'd870: toneL = `d;     15'd871: toneL = `d;
15'd872: toneL = `a;     15'd873: toneL = `a;
15'd874: toneL = `a;     15'd875: toneL = `a;
15'd876: toneL = `a;     15'd877: toneL = `a;
15'd878: toneL = `a;     15'd879: toneL = `a;
15'd880: toneL = `hd;     15'd881: toneL = `hd;
15'd882: toneL = `hd;     15'd883: toneL = `hd;
15'd884: toneL = `hd;     15'd885: toneL = `hd;
15'd886: toneL = `hd;     15'd887: toneL = `hd;
15'd888: toneL = `hd;     15'd889: toneL = `hd;
15'd890: toneL = `hd;     15'd891: toneL = `hd;
15'd892: toneL = `hd;     15'd893: toneL = `hd;
15'd894: toneL = `hd;     15'd895: toneL = `hd;
15'd896: toneL = `e;     15'd897: toneL = `e;
15'd898: toneL = `e;     15'd899: toneL = `e;
15'd900: toneL = `e;     15'd901: toneL = `e;
15'd902: toneL = `e;     15'd903: toneL = `e;
15'd904: toneL = `b;     15'd905: toneL = `b;
15'd906: toneL = `b;     15'd907: toneL = `b;
15'd908: toneL = `b;     15'd909: toneL = `b;
15'd910: toneL = `b;     15'd911: toneL = `b;
15'd912: toneL = `he;     15'd913: toneL = `he;
15'd914: toneL = `he;     15'd915: toneL = `he;
15'd916: toneL = `he;     15'd917: toneL = `he;
15'd918: toneL = `he;     15'd919: toneL = `he;
15'd920: toneL = `he;     15'd921: toneL = `he;
15'd922: toneL = `he;     15'd923: toneL = `he;
15'd924: toneL = `he;     15'd925: toneL = `he;
15'd926: toneL = `he;     15'd927: toneL = `he;
15'd928: toneL = `a;     15'd929: toneL = `a;
15'd930: toneL = `a;     15'd931: toneL = `a;
15'd932: toneL = `a;     15'd933: toneL = `a;
15'd934: toneL = `a;     15'd935: toneL = `a;
15'd936: toneL = `he;     15'd937: toneL = `he;
15'd938: toneL = `he;     15'd939: toneL = `he;
15'd940: toneL = `he;     15'd941: toneL = `he;
15'd942: toneL = `he;     15'd943: toneL = `he;
15'd944: toneL = `ha;     15'd945: toneL = `ha;
15'd946: toneL = `ha;     15'd947: toneL = `ha;
15'd948: toneL = `ha;     15'd949: toneL = `ha;
15'd950: toneL = `ha;     15'd951: toneL = `ha;
15'd952: toneL = `ha;     15'd953: toneL = `ha;
15'd954: toneL = `ha;     15'd955: toneL = `ha;
15'd956: toneL = `ha;     15'd957: toneL = `ha;
15'd958: toneL = `ha;     15'd959: toneL = `ha;
15'd960: toneL = `f;     15'd961: toneL = `f;
15'd962: toneL = `f;     15'd963: toneL = `f;
15'd964: toneL = `f;     15'd965: toneL = `f;
15'd966: toneL = `f;     15'd967: toneL = `f;
15'd968: toneL = `hc;     15'd969: toneL = `hc;
15'd970: toneL = `hc;     15'd971: toneL = `hc;
15'd972: toneL = `hc;     15'd973: toneL = `hc;
15'd974: toneL = `hc;     15'd975: toneL = `hc;
15'd976: toneL = `hf;     15'd977: toneL = `hf;
15'd978: toneL = `hf;     15'd979: toneL = `hf;
15'd980: toneL = `hf;     15'd981: toneL = `hf;
15'd982: toneL = `hf;     15'd983: toneL = `hf;
15'd984: toneL = `hf;     15'd985: toneL = `hf;
15'd986: toneL = `hf;     15'd987: toneL = `hf;
15'd988: toneL = `hf;     15'd989: toneL = `hf;
15'd990: toneL = `hf;     15'd991: toneL = `hf;
15'd992: toneL = `e;     15'd993: toneL = `e;
15'd994: toneL = `e;     15'd995: toneL = `e;
15'd996: toneL = `e;     15'd997: toneL = `e;
15'd998: toneL = `e;     15'd999: toneL = `e;
15'd1000: toneL = `b;     15'd1001: toneL = `b;
15'd1002: toneL = `b;     15'd1003: toneL = `b;
15'd1004: toneL = `b;     15'd1005: toneL = `b;
15'd1006: toneL = `b;     15'd1007: toneL = `b;
15'd1008: toneL = `he;     15'd1009: toneL = `he;
15'd1010: toneL = `he;     15'd1011: toneL = `he;
15'd1012: toneL = `he;     15'd1013: toneL = `he;
15'd1014: toneL = `he;     15'd1015: toneL = `he;
15'd1016: toneL = `he;     15'd1017: toneL = `he;
15'd1018: toneL = `he;     15'd1019: toneL = `he;
15'd1020: toneL = `he;     15'd1021: toneL = `he;
15'd1022: toneL = `he;     15'd1023: toneL = `he;
15'd1024: toneL = `a;     15'd1025: toneL = `a;
15'd1026: toneL = `a;     15'd1027: toneL = `a;
15'd1028: toneL = `a;     15'd1029: toneL = `a;
15'd1030: toneL = `a;     15'd1031: toneL = `a;
15'd1032: toneL = `he;     15'd1033: toneL = `he;
15'd1034: toneL = `he;     15'd1035: toneL = `he;
15'd1036: toneL = `he;     15'd1037: toneL = `he;
15'd1038: toneL = `he;     15'd1039: toneL = `he;
15'd1040: toneL = `ha;     15'd1041: toneL = `ha;
15'd1042: toneL = `ha;     15'd1043: toneL = `ha;
15'd1044: toneL = `ha;     15'd1045: toneL = `ha;
15'd1046: toneL = `ha;     15'd1047: toneL = `ha;
15'd1048: toneL = `sil;     15'd1049: toneL = `ha;
15'd1050: toneL = `ha;     15'd1051: toneL = `ha;
15'd1052: toneL = `ha;     15'd1053: toneL = `ha;
15'd1054: toneL = `ha;     15'd1055: toneL = `ha;
15'd1056: toneL = `ha;     15'd1057: toneL = `ha;
15'd1058: toneL = `ha;     15'd1059: toneL = `ha;
15'd1060: toneL = `ha;     15'd1061: toneL = `ha;
15'd1062: toneL = `ha;     15'd1063: toneL = `ha;
15'd1064: toneL = `he;     15'd1065: toneL = `he;
15'd1066: toneL = `he;     15'd1067: toneL = `he;
15'd1068: toneL = `he;     15'd1069: toneL = `he;
15'd1070: toneL = `he;     15'd1071: toneL = `he;
15'd1072: toneL = `ha;     15'd1073: toneL = `ha;
15'd1074: toneL = `ha;     15'd1075: toneL = `ha;
15'd1076: toneL = `ha;     15'd1077: toneL = `ha;
15'd1078: toneL = `ha;     15'd1079: toneL = `ha;
15'd1080: toneL = `he;     15'd1081: toneL = `he;
15'd1082: toneL = `he;     15'd1083: toneL = `he;
15'd1084: toneL = `he;     15'd1085: toneL = `he;
15'd1086: toneL = `he;     15'd1087: toneL = `he;
15'd1088: toneL = `a;     15'd1089: toneL = `a;
15'd1090: toneL = `a;     15'd1091: toneL = `a;
15'd1092: toneL = `a;     15'd1093: toneL = `a;
15'd1094: toneL = `a;     15'd1095: toneL = `a;
15'd1096: toneL = `he;     15'd1097: toneL = `he;
15'd1098: toneL = `he;     15'd1099: toneL = `he;
15'd1100: toneL = `he;     15'd1101: toneL = `he;
15'd1102: toneL = `he;     15'd1103: toneL = `he;
15'd1104: toneL = `hb;     15'd1105: toneL = `hb;
15'd1106: toneL = `hb;     15'd1107: toneL = `hb;
15'd1108: toneL = `hb;     15'd1109: toneL = `hb;
15'd1110: toneL = `hb;     15'd1111: toneL = `hb;
15'd1112: toneL = `ha;     15'd1113: toneL = `ha;
15'd1114: toneL = `ha;     15'd1115: toneL = `ha;
15'd1116: toneL = `ha;     15'd1117: toneL = `ha;
15'd1118: toneL = `ha;     15'd1119: toneL = `ha;
15'd1120: toneL = `hhc;     15'd1121: toneL = `hhc;
15'd1122: toneL = `hhc;     15'd1123: toneL = `hhc;
15'd1124: toneL = `hhc;     15'd1125: toneL = `hhc;
15'd1126: toneL = `hhc;     15'd1127: toneL = `hhc;
15'd1128: toneL = `ha;     15'd1129: toneL = `ha;
15'd1130: toneL = `ha;     15'd1131: toneL = `ha;
15'd1132: toneL = `ha;     15'd1133: toneL = `ha;
15'd1134: toneL = `ha;     15'd1135: toneL = `ha;
15'd1136: toneL = `hb;     15'd1137: toneL = `hb;
15'd1138: toneL = `hb;     15'd1139: toneL = `hb;
15'd1140: toneL = `hb;     15'd1141: toneL = `hb;
15'd1142: toneL = `hb;     15'd1143: toneL = `hb;
15'd1144: toneL = `ha;     15'd1145: toneL = `ha;
15'd1146: toneL = `ha;     15'd1147: toneL = `ha;
15'd1148: toneL = `ha;     15'd1149: toneL = `ha;
15'd1150: toneL = `ha;     15'd1151: toneL = `ha;
15'd1152: toneL = `d;     15'd1153: toneL = `d;
15'd1154: toneL = `d;     15'd1155: toneL = `d;
15'd1156: toneL = `d;     15'd1157: toneL = `d;
15'd1158: toneL = `d;     15'd1159: toneL = `d;
15'd1160: toneL = `a;     15'd1161: toneL = `a;
15'd1162: toneL = `a;     15'd1163: toneL = `a;
15'd1164: toneL = `a;     15'd1165: toneL = `a;
15'd1166: toneL = `a;     15'd1167: toneL = `a;
15'd1168: toneL = `hd;     15'd1169: toneL = `hd;
15'd1170: toneL = `hd;     15'd1171: toneL = `hd;
15'd1172: toneL = `hd;     15'd1173: toneL = `hd;
15'd1174: toneL = `hd;     15'd1175: toneL = `hd;
15'd1176: toneL = `a;     15'd1177: toneL = `a;
15'd1178: toneL = `a;     15'd1179: toneL = `a;
15'd1180: toneL = `a;     15'd1181: toneL = `a;
15'd1182: toneL = `a;     15'd1183: toneL = `a;
15'd1184: toneL = `e;     15'd1185: toneL = `e;
15'd1186: toneL = `e;     15'd1187: toneL = `e;
15'd1188: toneL = `e;     15'd1189: toneL = `e;
15'd1190: toneL = `e;     15'd1191: toneL = `e;
15'd1192: toneL = `b;     15'd1193: toneL = `b;
15'd1194: toneL = `b;     15'd1195: toneL = `b;
15'd1196: toneL = `b;     15'd1197: toneL = `b;
15'd1198: toneL = `b;     15'd1199: toneL = `b;
15'd1200: toneL = `he;     15'd1201: toneL = `he;
15'd1202: toneL = `he;     15'd1203: toneL = `he;
15'd1204: toneL = `he;     15'd1205: toneL = `he;
15'd1206: toneL = `he;     15'd1207: toneL = `he;
15'd1208: toneL = `b;     15'd1209: toneL = `b;
15'd1210: toneL = `b;     15'd1211: toneL = `b;
15'd1212: toneL = `b;     15'd1213: toneL = `b;
15'd1214: toneL = `b;     15'd1215: toneL = `b;
                    default: toneL = `sil;
                endcase
            end
            else begin
                case(ibeatNum)
                    15'd0: toneL = `hc;     15'd1: toneL = `hc;
                    15'd2: toneL = `hc;     15'd3: toneL = `hc;
                    15'd4: toneL = `hc;     15'd5: toneL = `hc;
                    15'd6: toneL = `hc;     15'd7: toneL = `hc;
                    15'd8: toneL = `hc;     15'd9: toneL = `hc;
                    15'd10: toneL = `hc;     15'd11: toneL = `hc;
                    15'd12: toneL = `hc;     15'd13: toneL = `hc;
                    15'd14: toneL = `hc;     15'd15: toneL = `hc;
                    15'd16: toneL = `hc;     15'd17: toneL = `hc;
                    15'd18: toneL = `hc;     15'd19: toneL = `hc;
                    15'd20: toneL = `hc;     15'd21: toneL = `hc;
                    15'd22: toneL = `hc;     15'd23: toneL = `hc;
                    15'd24: toneL = `hc;     15'd25: toneL = `hc;
                    15'd26: toneL = `hc;     15'd27: toneL = `hc;
                    15'd28: toneL = `hc;     15'd29: toneL = `hc;
                    15'd30: toneL = `hc;     15'd31: toneL = `hc;
                    15'd32: toneL = `g;     15'd33: toneL = `g;
                    15'd34: toneL = `g;     15'd35: toneL = `g;
                    15'd36: toneL = `g;     15'd37: toneL = `g;
                    15'd38: toneL = `g;     15'd39: toneL = `g;
                    15'd40: toneL = `g;     15'd41: toneL = `g;
                    15'd42: toneL = `g;     15'd43: toneL = `g;
                    15'd44: toneL = `g;     15'd45: toneL = `g;
                    15'd46: toneL = `g;     15'd47: toneL = `g;
                    15'd48: toneL = `g;     15'd49: toneL = `g;
                    15'd50: toneL = `g;     15'd51: toneL = `g;
                    15'd52: toneL = `g;     15'd53: toneL = `g;
                    15'd54: toneL = `g;     15'd55: toneL = `g;
                    15'd56: toneL = `g;     15'd57: toneL = `g;
                    15'd58: toneL = `g;     15'd59: toneL = `g;
                    15'd60: toneL = `g;     15'd61: toneL = `g;
                    15'd62: toneL = `g;     15'd63: toneL = `g;
                    15'd64: toneL = `hc;     15'd65: toneL = `hc;
                    15'd66: toneL = `hc;     15'd67: toneL = `hc;
                    15'd68: toneL = `hc;     15'd69: toneL = `hc;
                    15'd70: toneL = `hc;     15'd71: toneL = `hc;
                    15'd72: toneL = `hc;     15'd73: toneL = `hc;
                    15'd74: toneL = `hc;     15'd75: toneL = `hc;
                    15'd76: toneL = `hc;     15'd77: toneL = `hc;
                    15'd78: toneL = `hc;     15'd79: toneL = `hc;
                    15'd80: toneL = `hc;     15'd81: toneL = `hc;
                    15'd82: toneL = `hc;     15'd83: toneL = `hc;
                    15'd84: toneL = `hc;     15'd85: toneL = `hc;
                    15'd86: toneL = `hc;     15'd87: toneL = `hc;
                    15'd88: toneL = `hc;     15'd89: toneL = `hc;
                    15'd90: toneL = `hc;     15'd91: toneL = `hc;
                    15'd92: toneL = `hc;     15'd93: toneL = `hc;
                    15'd94: toneL = `hc;     15'd95: toneL = `hc;
                    15'd96: toneL = `g;     15'd97: toneL = `g;
                    15'd98: toneL = `g;     15'd99: toneL = `g;
                    15'd100: toneL = `g;     15'd101: toneL = `g;
                    15'd102: toneL = `g;     15'd103: toneL = `g;
                    15'd104: toneL = `g;     15'd105: toneL = `g;
                    15'd106: toneL = `g;     15'd107: toneL = `g;
                    15'd108: toneL = `g;     15'd109: toneL = `g;
                    15'd110: toneL = `g;     15'd111: toneL = `g;
                    15'd112: toneL = `g;     15'd113: toneL = `g;
                    15'd114: toneL = `g;     15'd115: toneL = `g;
                    15'd116: toneL = `g;     15'd117: toneL = `g;
                    15'd118: toneL = `g;     15'd119: toneL = `g;
                    15'd120: toneL = `g;     15'd121: toneL = `g;
                    15'd122: toneL = `g;     15'd123: toneL = `g;
                    15'd124: toneL = `g;     15'd125: toneL = `g;
                    15'd126: toneL = `g;     15'd127: toneL = `g;
                    15'd128: toneL = `c;     15'd129: toneL = `c;
                    15'd130: toneL = `c;     15'd131: toneL = `c;
                    15'd132: toneL = `c;     15'd133: toneL = `c;
                    15'd134: toneL = `c;     15'd135: toneL = `c;
                    15'd136: toneL = `c;     15'd137: toneL = `c;
                    15'd138: toneL = `c;     15'd139: toneL = `c;
                    15'd140: toneL = `c;     15'd141: toneL = `c;
                    15'd142: toneL = `c;     15'd143: toneL = `c;
                    15'd144: toneL = `d;     15'd145: toneL = `d;
                    15'd146: toneL = `d;     15'd147: toneL = `d;
                    15'd148: toneL = `d;     15'd149: toneL = `d;
                    15'd150: toneL = `d;     15'd151: toneL = `d;
                    15'd152: toneL = `d;     15'd153: toneL = `d;
                    15'd154: toneL = `d;     15'd155: toneL = `d;
                    15'd156: toneL = `d;     15'd157: toneL = `d;
                    15'd158: toneL = `d;     15'd159: toneL = `d;
                    15'd160: toneL = `e;     15'd161: toneL = `e;
                    15'd162: toneL = `e;     15'd163: toneL = `e;
                    15'd164: toneL = `e;     15'd165: toneL = `e;
                    15'd166: toneL = `e;     15'd167: toneL = `e;
                    15'd168: toneL = `e;     15'd169: toneL = `e;
                    15'd170: toneL = `e;     15'd171: toneL = `e;
                    15'd172: toneL = `e;     15'd173: toneL = `e;
                    15'd174: toneL = `e;     15'd175: toneL = `e;
                    15'd176: toneL = `e;     15'd177: toneL = `e;
                    15'd178: toneL = `e;     15'd179: toneL = `e;
                    15'd180: toneL = `e;     15'd181: toneL = `e;
                    15'd182: toneL = `e;     15'd183: toneL = `e;
                    15'd184: toneL = `e;     15'd185: toneL = `e;
                    15'd186: toneL = `e;     15'd187: toneL = `e;
                    15'd188: toneL = `e;     15'd189: toneL = `e;
                    15'd190: toneL = `e;     15'd191: toneL = `e;
                    15'd192: toneL = `c;     15'd193: toneL = `c;
                    15'd194: toneL = `c;     15'd195: toneL = `c;
                    15'd196: toneL = `c;     15'd197: toneL = `c;
                    15'd198: toneL = `c;     15'd199: toneL = `c;
                    15'd200: toneL = `c;     15'd201: toneL = `c;
                    15'd202: toneL = `c;     15'd203: toneL = `c;
                    15'd204: toneL = `c;     15'd205: toneL = `c;
                    15'd206: toneL = `c;     15'd207: toneL = `c;
                    15'd208: toneL = `d;     15'd209: toneL = `d;
                    15'd210: toneL = `d;     15'd211: toneL = `d;
                    15'd212: toneL = `d;     15'd213: toneL = `d;
                    15'd214: toneL = `d;     15'd215: toneL = `d;
                    15'd216: toneL = `d;     15'd217: toneL = `d;
                    15'd218: toneL = `d;     15'd219: toneL = `d;
                    15'd220: toneL = `d;     15'd221: toneL = `d;
                    15'd222: toneL = `d;     15'd223: toneL = `d;
                    15'd224: toneL = `e;     15'd225: toneL = `e;
                    15'd226: toneL = `e;     15'd227: toneL = `e;
                    15'd228: toneL = `e;     15'd229: toneL = `e;
                    15'd230: toneL = `e;     15'd231: toneL = `e;
                    15'd232: toneL = `e;     15'd233: toneL = `e;
                    15'd234: toneL = `e;     15'd235: toneL = `e;
                    15'd236: toneL = `e;     15'd237: toneL = `e;
                    15'd238: toneL = `e;     15'd239: toneL = `e;
                    15'd240: toneL = `e;     15'd241: toneL = `e;
                    15'd242: toneL = `e;     15'd243: toneL = `e;
                    15'd244: toneL = `e;     15'd245: toneL = `e;
                    15'd246: toneL = `e;     15'd247: toneL = `e;
                    15'd248: toneL = `e;     15'd249: toneL = `e;
                    15'd250: toneL = `e;     15'd251: toneL = `e;
                    15'd252: toneL = `e;     15'd253: toneL = `e;
                    15'd254: toneL = `e;     15'd255: toneL = `e;
                    15'd256: toneL = `e;     15'd257: toneL = `e;
                    15'd258: toneL = `e;     15'd259: toneL = `e;
                    15'd260: toneL = `e;     15'd261: toneL = `e;
                    15'd262: toneL = `e;     15'd263: toneL = `e;
                    15'd264: toneL = `e;     15'd265: toneL = `e;
                    15'd266: toneL = `e;     15'd267: toneL = `e;
                    15'd268: toneL = `e;     15'd269: toneL = `e;
                    15'd270: toneL = `e;     15'd271: toneL = `e;
                    15'd272: toneL = `f;     15'd273: toneL = `f;
                    15'd274: toneL = `f;     15'd275: toneL = `f;
                    15'd276: toneL = `f;     15'd277: toneL = `f;
                    15'd278: toneL = `f;     15'd279: toneL = `f;
                    15'd280: toneL = `f;     15'd281: toneL = `f;
                    15'd282: toneL = `f;     15'd283: toneL = `f;
                    15'd284: toneL = `f;     15'd285: toneL = `f;
                    15'd286: toneL = `f;     15'd287: toneL = `f;
                    15'd288: toneL = `g;     15'd289: toneL = `g;
                    15'd290: toneL = `g;     15'd291: toneL = `g;
                    15'd292: toneL = `g;     15'd293: toneL = `g;
                    15'd294: toneL = `g;     15'd295: toneL = `g;
                    15'd296: toneL = `g;     15'd297: toneL = `g;
                    15'd298: toneL = `g;     15'd299: toneL = `g;
                    15'd300: toneL = `g;     15'd301: toneL = `g;
                    15'd302: toneL = `g;     15'd303: toneL = `g;
                    15'd304: toneL = `g;     15'd305: toneL = `g;
                    15'd306: toneL = `g;     15'd307: toneL = `g;
                    15'd308: toneL = `g;     15'd309: toneL = `g;
                    15'd310: toneL = `g;     15'd311: toneL = `g;
                    15'd312: toneL = `g;     15'd313: toneL = `g;
                    15'd314: toneL = `g;     15'd315: toneL = `g;
                    15'd316: toneL = `g;     15'd317: toneL = `g;
                    15'd318: toneL = `g;     15'd319: toneL = `g;
                    15'd320: toneL = `e;     15'd321: toneL = `e;
                    15'd322: toneL = `e;     15'd323: toneL = `e;
                    15'd324: toneL = `e;     15'd325: toneL = `e;
                    15'd326: toneL = `e;     15'd327: toneL = `e;
                    15'd328: toneL = `e;     15'd329: toneL = `e;
                    15'd330: toneL = `e;     15'd331: toneL = `e;
                    15'd332: toneL = `e;     15'd333: toneL = `e;
                    15'd334: toneL = `e;     15'd335: toneL = `e;
                    15'd336: toneL = `f;     15'd337: toneL = `f;
                    15'd338: toneL = `f;     15'd339: toneL = `f;
                    15'd340: toneL = `f;     15'd341: toneL = `f;
                    15'd342: toneL = `f;     15'd343: toneL = `f;
                    15'd344: toneL = `f;     15'd345: toneL = `f;
                    15'd346: toneL = `f;     15'd347: toneL = `f;
                    15'd348: toneL = `f;     15'd349: toneL = `f;
                    15'd350: toneL = `f;     15'd351: toneL = `f;
                    15'd352: toneL = `g;     15'd353: toneL = `g;
                    15'd354: toneL = `g;     15'd355: toneL = `g;
                    15'd356: toneL = `g;     15'd357: toneL = `g;
                    15'd358: toneL = `g;     15'd359: toneL = `g;
                    15'd360: toneL = `g;     15'd361: toneL = `g;
                    15'd362: toneL = `g;     15'd363: toneL = `g;
                    15'd364: toneL = `g;     15'd365: toneL = `g;
                    15'd366: toneL = `g;     15'd367: toneL = `g;
                    15'd368: toneL = `g;     15'd369: toneL = `g;
                    15'd370: toneL = `g;     15'd371: toneL = `g;
                    15'd372: toneL = `g;     15'd373: toneL = `g;
                    15'd374: toneL = `g;     15'd375: toneL = `g;
                    15'd376: toneL = `sil;     15'd377: toneL = `sil;
                    15'd378: toneL = `g;     15'd379: toneL = `g;
                    15'd380: toneL = `g;     15'd381: toneL = `g;
                    15'd382: toneL = `g;     15'd383: toneL = `g;
                    15'd384: toneL = `g;     15'd385: toneL = `g;
                    15'd386: toneL = `g;     15'd387: toneL = `g;
                    15'd388: toneL = `g;     15'd389: toneL = `g;
                    15'd390: toneL = `g;     15'd391: toneL = `g;
                    15'd392: toneL = `g;     15'd393: toneL = `g;
                    15'd394: toneL = `g;     15'd395: toneL = `g;
                    15'd396: toneL = `g;     15'd397: toneL = `g;
                    15'd398: toneL = `g;     15'd399: toneL = `g;
                    15'd400: toneL = `g;     15'd401: toneL = `g;
                    15'd402: toneL = `g;     15'd403: toneL = `g;
                    15'd404: toneL = `g;     15'd405: toneL = `g;
                    15'd406: toneL = `g;     15'd407: toneL = `g;
                    15'd408: toneL = `g;     15'd409: toneL = `g;
                    15'd410: toneL = `g;     15'd411: toneL = `g;
                    15'd412: toneL = `g;     15'd413: toneL = `g;
                    15'd414: toneL = `g;     15'd415: toneL = `g;
                    15'd416: toneL = `e;     15'd417: toneL = `e;
                    15'd418: toneL = `e;     15'd419: toneL = `e;
                    15'd420: toneL = `e;     15'd421: toneL = `e;
                    15'd422: toneL = `e;     15'd423: toneL = `e;
                    15'd424: toneL = `e;     15'd425: toneL = `e;
                    15'd426: toneL = `e;     15'd427: toneL = `e;
                    15'd428: toneL = `e;     15'd429: toneL = `e;
                    15'd430: toneL = `e;     15'd431: toneL = `e;
                    15'd432: toneL = `e;     15'd433: toneL = `e;
                    15'd434: toneL = `e;     15'd435: toneL = `e;
                    15'd436: toneL = `e;     15'd437: toneL = `e;
                    15'd438: toneL = `e;     15'd439: toneL = `e;
                    15'd440: toneL = `e;     15'd441: toneL = `e;
                    15'd442: toneL = `e;     15'd443: toneL = `e;
                    15'd444: toneL = `e;     15'd445: toneL = `e;
                    15'd446: toneL = `e;     15'd447: toneL = `e;
                    15'd448: toneL = `g;     15'd449: toneL = `g;
                    15'd450: toneL = `g;     15'd451: toneL = `g;
                    15'd452: toneL = `g;     15'd453: toneL = `g;
                    15'd454: toneL = `g;     15'd455: toneL = `g;
                    15'd456: toneL = `g;     15'd457: toneL = `g;
                    15'd458: toneL = `g;     15'd459: toneL = `g;
                    15'd460: toneL = `g;     15'd461: toneL = `g;
                    15'd462: toneL = `g;     15'd463: toneL = `g;
                    15'd464: toneL = `g;     15'd465: toneL = `g;
                    15'd466: toneL = `g;     15'd467: toneL = `g;
                    15'd468: toneL = `g;     15'd469: toneL = `g;
                    15'd470: toneL = `g;     15'd471: toneL = `g;
                    15'd472: toneL = `g;     15'd473: toneL = `g;
                    15'd474: toneL = `g;     15'd475: toneL = `g;
                    15'd476: toneL = `g;     15'd477: toneL = `g;
                    15'd478: toneL = `g;     15'd479: toneL = `g;
                    15'd480: toneL = `e;     15'd481: toneL = `e;
                    15'd482: toneL = `e;     15'd483: toneL = `e;
                    15'd484: toneL = `e;     15'd485: toneL = `e;
                    15'd486: toneL = `e;     15'd487: toneL = `e;
                    15'd488: toneL = `e;     15'd489: toneL = `e;
                    15'd490: toneL = `e;     15'd491: toneL = `e;
                    15'd492: toneL = `e;     15'd493: toneL = `e;
                    15'd494: toneL = `e;     15'd495: toneL = `e;
                    15'd496: toneL = `e;     15'd497: toneL = `e;
                    15'd498: toneL = `e;     15'd499: toneL = `e;
                    15'd500: toneL = `e;     15'd501: toneL = `e;
                    15'd502: toneL = `e;     15'd503: toneL = `e;
                    15'd504: toneL = `e;     15'd505: toneL = `e;
                    15'd506: toneL = `e;     15'd507: toneL = `e;
                    15'd508: toneL = `e;     15'd509: toneL = `e;
                    15'd510: toneL = `e;     15'd511: toneL = `e;
                    default: toneL = `sil;
                endcase
            end
            //case(ibeatNum)
                // 12'd0: toneL = `hc;  	12'd1: toneL = `hc; // HC (two-beat)
                // 12'd2: toneL = `hc;  	12'd3: toneL = `hc;
                // 12'd4: toneL = `hc;	    12'd5: toneL = `hc;
                // 12'd6: toneL = `hc;  	12'd7: toneL = `hc;
                // 12'd8: toneL = `hc;	    12'd9: toneL = `hc;
                // 12'd10: toneL = `hc;	12'd11: toneL = `hc;
                // 12'd12: toneL = `hc;	12'd13: toneL = `hc;
                // 12'd14: toneL = `hc;	12'd15: toneL = `hc;

                // 12'd16: toneL = `hc;	12'd17: toneL = `hc;
                // 12'd18: toneL = `hc;	12'd19: toneL = `hc;
                // 12'd20: toneL = `hc;	12'd21: toneL = `hc;
                // 12'd22: toneL = `hc;	12'd23: toneL = `hc;
                // 12'd24: toneL = `hc;	12'd25: toneL = `hc;
                // 12'd26: toneL = `hc;	12'd27: toneL = `hc;
                // 12'd28: toneL = `hc;	12'd29: toneL = `hc;
                // 12'd30: toneL = `hc;	12'd31: toneL = `hc;

                // 12'd32: toneL = `g;	    12'd33: toneL = `g; // G (one-beat)
                // 12'd34: toneL = `g;	    12'd35: toneL = `g;
                // 12'd36: toneL = `g;	    12'd37: toneL = `g;
                // 12'd38: toneL = `g;	    12'd39: toneL = `g;
                // 12'd40: toneL = `g;	    12'd41: toneL = `g;
                // 12'd42: toneL = `g;	    12'd43: toneL = `g;
                // 12'd44: toneL = `g;	    12'd45: toneL = `g;
                // 12'd46: toneL = `g;	    12'd47: toneL = `g;

                // 12'd48: toneL = `b;	    12'd49: toneL = `b; // B (one-beat)
                // 12'd50: toneL = `b;	    12'd51: toneL = `b;
                // 12'd52: toneL = `b;	    12'd53: toneL = `b;
                // 12'd54: toneL = `b;	    12'd55: toneL = `b;
                // 12'd56: toneL = `b;	    12'd57: toneL = `b;
                // 12'd58: toneL = `b;	    12'd59: toneL = `b;
                // 12'd60: toneL = `b;	    12'd61: toneL = `b;
                // 12'd62: toneL = `b;	    12'd63: toneL = `b;

                // 12'd64: toneL = `hc;	    12'd65: toneL = `hc; // HC (two-beat)
                // 12'd66: toneL = `hc;	    12'd67: toneL = `hc;
                // 12'd68: toneL = `hc;	    12'd69: toneL = `hc;
                // 12'd70: toneL = `hc;	    12'd71: toneL = `hc;
                // 12'd72: toneL = `hc;	    12'd73: toneL = `hc;
                // 12'd74: toneL = `hc;	    12'd75: toneL = `hc;
                // 12'd76: toneL = `hc;	    12'd77: toneL = `hc;
                // 12'd78: toneL = `hc;	    12'd79: toneL = `hc;

                // 12'd80: toneL = `hc;	    12'd81: toneL = `hc;
                // 12'd82: toneL = `hc;	    12'd83: toneL = `hc;
                // 12'd84: toneL = `hc;	    12'd85: toneL = `hc;
                // 12'd86: toneL = `hc;	    12'd87: toneL = `hc;
                // 12'd88: toneL = `hc;	    12'd89: toneL = `hc;
                // 12'd90: toneL = `hc;	    12'd91: toneL = `hc;
                // 12'd92: toneL = `hc;	    12'd93: toneL = `hc;
                // 12'd94: toneL = `hc;	    12'd95: toneL = `hc;

                // 12'd96: toneL = `g;	    12'd97: toneL = `g; // G (one-beat)
                // 12'd98: toneL = `g; 	12'd99: toneL = `g;
                // 12'd100: toneL = `g;	12'd101: toneL = `g;
                // 12'd102: toneL = `g;	12'd103: toneL = `g;
                // 12'd104: toneL = `g;	12'd105: toneL = `g;
                // 12'd106: toneL = `g;	12'd107: toneL = `g;
                // 12'd108: toneL = `g;	12'd109: toneL = `g;
                // 12'd110: toneL = `g;	12'd111: toneL = `g;

                // 12'd112: toneL = `b;	12'd113: toneL = `b; // B (one-beat)
                // 12'd114: toneL = `b;	12'd115: toneL = `b;
                // 12'd116: toneL = `b;	12'd117: toneL = `b;
                // 12'd118: toneL = `b;	12'd119: toneL = `b;
                // 12'd120: toneL = `b;	12'd121: toneL = `b;
                // 12'd122: toneL = `b;	12'd123: toneL = `b;
                // 12'd124: toneL = `b;	12'd125: toneL = `b;
                // 12'd126: toneL = `b;	12'd127: toneL = `b;
                // 15'd0: toneL = `hd;     15'd1: toneL = `hd;
                //     15'd2: toneL = `hd;     15'd3: toneL = `hd;
                //     15'd4: toneL = `hd;     15'd5: toneL = `hd;
                //     15'd6: toneL = `hd;     15'd7: toneL = `hd;
                //     15'd8: toneL = `hd;     15'd9: toneL = `hd;
                //     15'd10: toneL = `hd;     15'd11: toneL = `hd;
                //     15'd12: toneL = `hd;     15'd13: toneL = `hd;
                //     15'd14: toneL = `hd;     15'd15: toneL = `hd;
                //     15'd16: toneL = `hd;     15'd17: toneL = `hd;
                //     15'd18: toneL = `hd;     15'd19: toneL = `hd;
                //     15'd20: toneL = `hd;     15'd21: toneL = `hd;
                //     15'd22: toneL = `hd;     15'd23: toneL = `hd;
                //     15'd24: toneL = `hd;     15'd25: toneL = `hd;
                //     15'd26: toneL = `hd;     15'd27: toneL = `hd;
                //     15'd28: toneL = `hd;     15'd29: toneL = `hd;
                //     15'd30: toneL = `hd;     15'd31: toneL = `hd;
                //     15'd32: toneL = `a;     15'd33: toneL = `a;
                //     15'd34: toneL = `a;     15'd35: toneL = `a;
                //     15'd36: toneL = `a;     15'd37: toneL = `a;
                //     15'd38: toneL = `a;     15'd39: toneL = `a;
                //     15'd40: toneL = `a;     15'd41: toneL = `a;
                //     15'd42: toneL = `a;     15'd43: toneL = `a;
                //     15'd44: toneL = `a;     15'd45: toneL = `a;
                //     15'd46: toneL = `a;     15'd47: toneL = `a;
                //     15'd48: toneL = `a;     15'd49: toneL = `a;
                //     15'd50: toneL = `a;     15'd51: toneL = `a;
                //     15'd52: toneL = `a;     15'd53: toneL = `a;
                //     15'd54: toneL = `a;     15'd55: toneL = `a;
                //     15'd56: toneL = `a;     15'd57: toneL = `a;
                //     15'd58: toneL = `a;     15'd59: toneL = `a;
                //     15'd60: toneL = `a;     15'd61: toneL = `a;
                //     15'd62: toneL = `a;     15'd63: toneL = `a;
                //     15'd64: toneL = `b;     15'd65: toneL = `b;
                //     15'd66: toneL = `b;     15'd67: toneL = `b;
                //     15'd68: toneL = `b;     15'd69: toneL = `b;
                //     15'd70: toneL = `b;     15'd71: toneL = `b;
                //     15'd72: toneL = `b;     15'd73: toneL = `b;
                //     15'd74: toneL = `b;     15'd75: toneL = `b;
                //     15'd76: toneL = `b;     15'd77: toneL = `b;
                //     15'd78: toneL = `b;     15'd79: toneL = `b;
                //     15'd80: toneL = `b;     15'd81: toneL = `b;
                //     15'd82: toneL = `b;     15'd83: toneL = `b;
                //     15'd84: toneL = `b;     15'd85: toneL = `b;
                //     15'd86: toneL = `b;     15'd87: toneL = `b;
                //     15'd88: toneL = `b;     15'd89: toneL = `b;
                //     15'd90: toneL = `b;     15'd91: toneL = `b;
                //     15'd92: toneL = `b;     15'd93: toneL = `b;
                //     15'd94: toneL = `b;     15'd95: toneL = `b;
                //     15'd96: toneL = `rf;     15'd97: toneL = `rf;
                //     15'd98: toneL = `rf;     15'd99: toneL = `rf;
                //     15'd100: toneL = `rf;     15'd101: toneL = `rf;
                //     15'd102: toneL = `rf;     15'd103: toneL = `rf;
                //     15'd104: toneL = `rf;     15'd105: toneL = `rf;
                //     15'd106: toneL = `rf;     15'd107: toneL = `rf;
                //     15'd108: toneL = `rf;     15'd109: toneL = `rf;
                //     15'd110: toneL = `rf;     15'd111: toneL = `rf;
                //     15'd112: toneL = `rf;     15'd113: toneL = `rf;
                //     15'd114: toneL = `rf;     15'd115: toneL = `rf;
                //     15'd116: toneL = `rf;     15'd117: toneL = `rf;
                //     15'd118: toneL = `rf;     15'd119: toneL = `rf;
                //     15'd120: toneL = `rf;     15'd121: toneL = `rf;
                //     15'd122: toneL = `rf;     15'd123: toneL = `rf;
                //     15'd124: toneL = `rf;     15'd125: toneL = `rf;
                //     15'd126: toneL = `rf;     15'd127: toneL = `rf;
                //     15'd128: toneL = `g;     15'd129: toneL = `g;
                //     15'd130: toneL = `g;     15'd131: toneL = `g;
                //     15'd132: toneL = `g;     15'd133: toneL = `g;
                //     15'd134: toneL = `g;     15'd135: toneL = `g;
                //     15'd136: toneL = `g;     15'd137: toneL = `g;
                //     15'd138: toneL = `g;     15'd139: toneL = `g;
                //     15'd140: toneL = `g;     15'd141: toneL = `g;
                //     15'd142: toneL = `g;     15'd143: toneL = `g;
                //     15'd144: toneL = `g;     15'd145: toneL = `g;
                //     15'd146: toneL = `g;     15'd147: toneL = `g;
                //     15'd148: toneL = `g;     15'd149: toneL = `g;
                //     15'd150: toneL = `g;     15'd151: toneL = `g;
                //     15'd152: toneL = `g;     15'd153: toneL = `g;
                //     15'd154: toneL = `g;     15'd155: toneL = `g;
                //     15'd156: toneL = `g;     15'd157: toneL = `g;
                //     15'd158: toneL = `g;     15'd159: toneL = `g;
                //     15'd160: toneL = `d;     15'd161: toneL = `d;
                //     15'd162: toneL = `d;     15'd163: toneL = `d;
                //     15'd164: toneL = `d;     15'd165: toneL = `d;
                //     15'd166: toneL = `d;     15'd167: toneL = `d;
                //     15'd168: toneL = `d;     15'd169: toneL = `d;
                //     15'd170: toneL = `d;     15'd171: toneL = `d;
                //     15'd172: toneL = `d;     15'd173: toneL = `d;
                //     15'd174: toneL = `d;     15'd175: toneL = `d;
                //     15'd176: toneL = `d;     15'd177: toneL = `d;
                //     15'd178: toneL = `d;     15'd179: toneL = `d;
                //     15'd180: toneL = `d;     15'd181: toneL = `d;
                //     15'd182: toneL = `d;     15'd183: toneL = `d;
                //     15'd184: toneL = `d;     15'd185: toneL = `d;
                //     15'd186: toneL = `d;     15'd187: toneL = `d;
                //     15'd188: toneL = `d;     15'd189: toneL = `d;
                //     15'd190: toneL = `d;     15'd191: toneL = `d;
                //     15'd192: toneL = `g;     15'd193: toneL = `g;
                //     15'd194: toneL = `g;     15'd195: toneL = `g;
                //     15'd196: toneL = `g;     15'd197: toneL = `g;
                //     15'd198: toneL = `g;     15'd199: toneL = `g;
                //     15'd200: toneL = `g;     15'd201: toneL = `g;
                //     15'd202: toneL = `g;     15'd203: toneL = `g;
                //     15'd204: toneL = `g;     15'd205: toneL = `g;
                //     15'd206: toneL = `g;     15'd207: toneL = `g;
                //     15'd208: toneL = `g;     15'd209: toneL = `g;
                //     15'd210: toneL = `g;     15'd211: toneL = `g;
                //     15'd212: toneL = `g;     15'd213: toneL = `g;
                //     15'd214: toneL = `g;     15'd215: toneL = `g;
                //     15'd216: toneL = `g;     15'd217: toneL = `g;
                //     15'd218: toneL = `g;     15'd219: toneL = `g;
                //     15'd220: toneL = `g;     15'd221: toneL = `g;
                //     15'd222: toneL = `g;     15'd223: toneL = `g;
                //     15'd224: toneL = `a;     15'd225: toneL = `a;
                //     15'd226: toneL = `a;     15'd227: toneL = `a;
                //     15'd228: toneL = `a;     15'd229: toneL = `a;
                //     15'd230: toneL = `a;     15'd231: toneL = `a;
                //     15'd232: toneL = `a;     15'd233: toneL = `a;
                //     15'd234: toneL = `a;     15'd235: toneL = `a;
                //     15'd236: toneL = `a;     15'd237: toneL = `a;
                //     15'd238: toneL = `a;     15'd239: toneL = `a;
                //     15'd240: toneL = `a;     15'd241: toneL = `a;
                //     15'd242: toneL = `a;     15'd243: toneL = `a;
                //     15'd244: toneL = `a;     15'd245: toneL = `a;
                //     15'd246: toneL = `a;     15'd247: toneL = `a;
                //     15'd248: toneL = `a;     15'd249: toneL = `a;
                //     15'd250: toneL = `a;     15'd251: toneL = `a;
                //     15'd252: toneL = `a;     15'd253: toneL = `a;
                //     15'd254: toneL = `a;     15'd255: toneL = `a;
                //     15'd256: toneL = `ha;     15'd257: toneL = `ha;
                //     15'd258: toneL = `ha;     15'd259: toneL = `ha;
                //     15'd260: toneL = `ha;     15'd261: toneL = `ha;
                //     15'd262: toneL = `ha;     15'd263: toneL = `ha;
                //     15'd264: toneL = `rhf;     15'd265: toneL = `rhf;
                //     15'd266: toneL = `rhf;     15'd267: toneL = `rhf;
                //     15'd268: toneL = `hg;     15'd269: toneL = `hg;
                //     15'd270: toneL = `hg;     15'd271: toneL = `hg;
                //     15'd272: toneL = `ha;     15'd273: toneL = `ha;
                //     15'd274: toneL = `ha;     15'd275: toneL = `ha;
                //     15'd276: toneL = `ha;     15'd277: toneL = `ha;
                //     15'd278: toneL = `ha;     15'd279: toneL = `ha;
                //     15'd280: toneL = `rhf;     15'd281: toneL = `rhf;
                //     15'd282: toneL = `rhf;     15'd283: toneL = `rhf;
                //     15'd284: toneL = `hg;     15'd285: toneL = `hg;
                //     15'd286: toneL = `hg;     15'd287: toneL = `hg;
                //     15'd288: toneL = `ha;     15'd289: toneL = `ha;
                //     15'd290: toneL = `ha;     15'd291: toneL = `ha;
                //     15'd292: toneL = `a;     15'd293: toneL = `a;
                //     15'd294: toneL = `a;     15'd295: toneL = `a;
                //     15'd296: toneL = `b;     15'd297: toneL = `b;
                //     15'd298: toneL = `b;     15'd299: toneL = `b;
                //     15'd300: toneL = `rhc;     15'd301: toneL = `rhc;
                //     15'd302: toneL = `rhc;     15'd303: toneL = `rhc;
                //     15'd304: toneL = `hd;     15'd305: toneL = `hd;
                //     15'd306: toneL = `hd;     15'd307: toneL = `hd;
                //     15'd308: toneL = `he;     15'd309: toneL = `he;
                //     15'd310: toneL = `he;     15'd311: toneL = `he;
                //     15'd312: toneL = `rhf;     15'd313: toneL = `rhf;
                //     15'd314: toneL = `rhf;     15'd315: toneL = `rhf;
                //     15'd316: toneL = `hg;     15'd317: toneL = `hg;
                //     15'd318: toneL = `hg;     15'd319: toneL = `hg;

                    // 15'd0: toneL = `hc;     15'd1: toneL = `hc;
                    // 15'd2: toneL = `hc;     15'd3: toneL = `hc;
                    // 15'd4: toneL = `hc;     15'd5: toneL = `hc;
                    // 15'd6: toneL = `hc;     15'd7: toneL = `hc;
                    // 15'd8: toneL = `hc;     15'd9: toneL = `hc;
                    // 15'd10: toneL = `hc;     15'd11: toneL = `hc;
                    // 15'd12: toneL = `hc;     15'd13: toneL = `hc;
                    // 15'd14: toneL = `hc;     15'd15: toneL = `hc;
                    // 15'd16: toneL = `hc;     15'd17: toneL = `hc;
                    // 15'd18: toneL = `hc;     15'd19: toneL = `hc;
                    // 15'd20: toneL = `hc;     15'd21: toneL = `hc;
                    // 15'd22: toneL = `hc;     15'd23: toneL = `hc;
                    // 15'd24: toneL = `hc;     15'd25: toneL = `hc;
                    // 15'd26: toneL = `hc;     15'd27: toneL = `hc;
                    // 15'd28: toneL = `hc;     15'd29: toneL = `hc;
                    // 15'd30: toneL = `hc;     15'd31: toneL = `hc;
                    // 15'd32: toneL = `g;     15'd33: toneL = `g;
                    // 15'd34: toneL = `g;     15'd35: toneL = `g;
                    // 15'd36: toneL = `g;     15'd37: toneL = `g;
                    // 15'd38: toneL = `g;     15'd39: toneL = `g;
                    // 15'd40: toneL = `g;     15'd41: toneL = `g;
                    // 15'd42: toneL = `g;     15'd43: toneL = `g;
                    // 15'd44: toneL = `g;     15'd45: toneL = `g;
                    // 15'd46: toneL = `g;     15'd47: toneL = `g;
                    // 15'd48: toneL = `g;     15'd49: toneL = `g;
                    // 15'd50: toneL = `g;     15'd51: toneL = `g;
                    // 15'd52: toneL = `g;     15'd53: toneL = `g;
                    // 15'd54: toneL = `g;     15'd55: toneL = `g;
                    // 15'd56: toneL = `g;     15'd57: toneL = `g;
                    // 15'd58: toneL = `g;     15'd59: toneL = `g;
                    // 15'd60: toneL = `g;     15'd61: toneL = `g;
                    // 15'd62: toneL = `g;     15'd63: toneL = `g;
                    // 15'd64: toneL = `hc;     15'd65: toneL = `hc;
                    // 15'd66: toneL = `hc;     15'd67: toneL = `hc;
                    // 15'd68: toneL = `hc;     15'd69: toneL = `hc;
                    // 15'd70: toneL = `hc;     15'd71: toneL = `hc;
                    // 15'd72: toneL = `hc;     15'd73: toneL = `hc;
                    // 15'd74: toneL = `hc;     15'd75: toneL = `hc;
                    // 15'd76: toneL = `hc;     15'd77: toneL = `hc;
                    // 15'd78: toneL = `hc;     15'd79: toneL = `hc;
                    // 15'd80: toneL = `hc;     15'd81: toneL = `hc;
                    // 15'd82: toneL = `hc;     15'd83: toneL = `hc;
                    // 15'd84: toneL = `hc;     15'd85: toneL = `hc;
                    // 15'd86: toneL = `hc;     15'd87: toneL = `hc;
                    // 15'd88: toneL = `hc;     15'd89: toneL = `hc;
                    // 15'd90: toneL = `hc;     15'd91: toneL = `hc;
                    // 15'd92: toneL = `hc;     15'd93: toneL = `hc;
                    // 15'd94: toneL = `hc;     15'd95: toneL = `hc;
                    // 15'd96: toneL = `g;     15'd97: toneL = `g;
                    // 15'd98: toneL = `g;     15'd99: toneL = `g;
                    // 15'd100: toneL = `g;     15'd101: toneL = `g;
                    // 15'd102: toneL = `g;     15'd103: toneL = `g;
                    // 15'd104: toneL = `g;     15'd105: toneL = `g;
                    // 15'd106: toneL = `g;     15'd107: toneL = `g;
                    // 15'd108: toneL = `g;     15'd109: toneL = `g;
                    // 15'd110: toneL = `g;     15'd111: toneL = `g;
                    // 15'd112: toneL = `g;     15'd113: toneL = `g;
                    // 15'd114: toneL = `g;     15'd115: toneL = `g;
                    // 15'd116: toneL = `g;     15'd117: toneL = `g;
                    // 15'd118: toneL = `g;     15'd119: toneL = `g;
                    // 15'd120: toneL = `g;     15'd121: toneL = `g;
                    // 15'd122: toneL = `g;     15'd123: toneL = `g;
                    // 15'd124: toneL = `g;     15'd125: toneL = `g;
                    // 15'd126: toneL = `g;     15'd127: toneL = `g;
                    // 15'd128: toneL = `c;     15'd129: toneL = `c;
                    // 15'd130: toneL = `c;     15'd131: toneL = `c;
                    // 15'd132: toneL = `c;     15'd133: toneL = `c;
                    // 15'd134: toneL = `c;     15'd135: toneL = `c;
                    // 15'd136: toneL = `c;     15'd137: toneL = `c;
                    // 15'd138: toneL = `c;     15'd139: toneL = `c;
                    // 15'd140: toneL = `c;     15'd141: toneL = `c;
                    // 15'd142: toneL = `c;     15'd143: toneL = `c;
                    // 15'd144: toneL = `d;     15'd145: toneL = `d;
                    // 15'd146: toneL = `d;     15'd147: toneL = `d;
                    // 15'd148: toneL = `d;     15'd149: toneL = `d;
                    // 15'd150: toneL = `d;     15'd151: toneL = `d;
                    // 15'd152: toneL = `d;     15'd153: toneL = `d;
                    // 15'd154: toneL = `d;     15'd155: toneL = `d;
                    // 15'd156: toneL = `d;     15'd157: toneL = `d;
                    // 15'd158: toneL = `d;     15'd159: toneL = `d;
                    // 15'd160: toneL = `e;     15'd161: toneL = `e;
                    // 15'd162: toneL = `e;     15'd163: toneL = `e;
                    // 15'd164: toneL = `e;     15'd165: toneL = `e;
                    // 15'd166: toneL = `e;     15'd167: toneL = `e;
                    // 15'd168: toneL = `e;     15'd169: toneL = `e;
                    // 15'd170: toneL = `e;     15'd171: toneL = `e;
                    // 15'd172: toneL = `e;     15'd173: toneL = `e;
                    // 15'd174: toneL = `e;     15'd175: toneL = `e;
                    // 15'd176: toneL = `e;     15'd177: toneL = `e;
                    // 15'd178: toneL = `e;     15'd179: toneL = `e;
                    // 15'd180: toneL = `e;     15'd181: toneL = `e;
                    // 15'd182: toneL = `e;     15'd183: toneL = `e;
                    // 15'd184: toneL = `e;     15'd185: toneL = `e;
                    // 15'd186: toneL = `e;     15'd187: toneL = `e;
                    // 15'd188: toneL = `e;     15'd189: toneL = `e;
                    // 15'd190: toneL = `e;     15'd191: toneL = `e;
                    // 15'd192: toneL = `c;     15'd193: toneL = `c;
                    // 15'd194: toneL = `c;     15'd195: toneL = `c;
                    // 15'd196: toneL = `c;     15'd197: toneL = `c;
                    // 15'd198: toneL = `c;     15'd199: toneL = `c;
                    // 15'd200: toneL = `c;     15'd201: toneL = `c;
                    // 15'd202: toneL = `c;     15'd203: toneL = `c;
                    // 15'd204: toneL = `c;     15'd205: toneL = `c;
                    // 15'd206: toneL = `c;     15'd207: toneL = `c;
                    // 15'd208: toneL = `d;     15'd209: toneL = `d;
                    // 15'd210: toneL = `d;     15'd211: toneL = `d;
                    // 15'd212: toneL = `d;     15'd213: toneL = `d;
                    // 15'd214: toneL = `d;     15'd215: toneL = `d;
                    // 15'd216: toneL = `d;     15'd217: toneL = `d;
                    // 15'd218: toneL = `d;     15'd219: toneL = `d;
                    // 15'd220: toneL = `d;     15'd221: toneL = `d;
                    // 15'd222: toneL = `d;     15'd223: toneL = `d;
                    // 15'd224: toneL = `e;     15'd225: toneL = `e;
                    // 15'd226: toneL = `e;     15'd227: toneL = `e;
                    // 15'd228: toneL = `e;     15'd229: toneL = `e;
                    // 15'd230: toneL = `e;     15'd231: toneL = `e;
                    // 15'd232: toneL = `e;     15'd233: toneL = `e;
                    // 15'd234: toneL = `e;     15'd235: toneL = `e;
                    // 15'd236: toneL = `e;     15'd237: toneL = `e;
                    // 15'd238: toneL = `e;     15'd239: toneL = `e;
                    // 15'd240: toneL = `e;     15'd241: toneL = `e;
                    // 15'd242: toneL = `e;     15'd243: toneL = `e;
                    // 15'd244: toneL = `e;     15'd245: toneL = `e;
                    // 15'd246: toneL = `e;     15'd247: toneL = `e;
                    // 15'd248: toneL = `e;     15'd249: toneL = `e;
                    // 15'd250: toneL = `e;     15'd251: toneL = `e;
                    // 15'd252: toneL = `e;     15'd253: toneL = `e;
                    // 15'd254: toneL = `e;     15'd255: toneL = `e;
                    // 15'd256: toneL = `e;     15'd257: toneL = `e;
                    // 15'd258: toneL = `e;     15'd259: toneL = `e;
                    // 15'd260: toneL = `e;     15'd261: toneL = `e;
                    // 15'd262: toneL = `e;     15'd263: toneL = `e;
                    // 15'd264: toneL = `e;     15'd265: toneL = `e;
                    // 15'd266: toneL = `e;     15'd267: toneL = `e;
                    // 15'd268: toneL = `e;     15'd269: toneL = `e;
                    // 15'd270: toneL = `e;     15'd271: toneL = `e;
                    // 15'd272: toneL = `f;     15'd273: toneL = `f;
                    // 15'd274: toneL = `f;     15'd275: toneL = `f;
                    // 15'd276: toneL = `f;     15'd277: toneL = `f;
                    // 15'd278: toneL = `f;     15'd279: toneL = `f;
                    // 15'd280: toneL = `f;     15'd281: toneL = `f;
                    // 15'd282: toneL = `f;     15'd283: toneL = `f;
                    // 15'd284: toneL = `f;     15'd285: toneL = `f;
                    // 15'd286: toneL = `f;     15'd287: toneL = `f;
                    // 15'd288: toneL = `g;     15'd289: toneL = `g;
                    // 15'd290: toneL = `g;     15'd291: toneL = `g;
                    // 15'd292: toneL = `g;     15'd293: toneL = `g;
                    // 15'd294: toneL = `g;     15'd295: toneL = `g;
                    // 15'd296: toneL = `g;     15'd297: toneL = `g;
                    // 15'd298: toneL = `g;     15'd299: toneL = `g;
                    // 15'd300: toneL = `g;     15'd301: toneL = `g;
                    // 15'd302: toneL = `g;     15'd303: toneL = `g;
                    // 15'd304: toneL = `g;     15'd305: toneL = `g;
                    // 15'd306: toneL = `g;     15'd307: toneL = `g;
                    // 15'd308: toneL = `g;     15'd309: toneL = `g;
                    // 15'd310: toneL = `g;     15'd311: toneL = `g;
                    // 15'd312: toneL = `g;     15'd313: toneL = `g;
                    // 15'd314: toneL = `g;     15'd315: toneL = `g;
                    // 15'd316: toneL = `g;     15'd317: toneL = `g;
                    // 15'd318: toneL = `g;     15'd319: toneL = `g;
                    // 15'd320: toneL = `e;     15'd321: toneL = `e;
                    // 15'd322: toneL = `e;     15'd323: toneL = `e;
                    // 15'd324: toneL = `e;     15'd325: toneL = `e;
                    // 15'd326: toneL = `e;     15'd327: toneL = `e;
                    // 15'd328: toneL = `e;     15'd329: toneL = `e;
                    // 15'd330: toneL = `e;     15'd331: toneL = `e;
                    // 15'd332: toneL = `e;     15'd333: toneL = `e;
                    // 15'd334: toneL = `e;     15'd335: toneL = `e;
                    // 15'd336: toneL = `f;     15'd337: toneL = `f;
                    // 15'd338: toneL = `f;     15'd339: toneL = `f;
                    // 15'd340: toneL = `f;     15'd341: toneL = `f;
                    // 15'd342: toneL = `f;     15'd343: toneL = `f;
                    // 15'd344: toneL = `f;     15'd345: toneL = `f;
                    // 15'd346: toneL = `f;     15'd347: toneL = `f;
                    // 15'd348: toneL = `f;     15'd349: toneL = `f;
                    // 15'd350: toneL = `f;     15'd351: toneL = `f;
                    // 15'd352: toneL = `g;     15'd353: toneL = `g;
                    // 15'd354: toneL = `g;     15'd355: toneL = `g;
                    // 15'd356: toneL = `g;     15'd357: toneL = `g;
                    // 15'd358: toneL = `g;     15'd359: toneL = `g;
                    // 15'd360: toneL = `g;     15'd361: toneL = `g;
                    // 15'd362: toneL = `g;     15'd363: toneL = `g;
                    // 15'd364: toneL = `g;     15'd365: toneL = `g;
                    // 15'd366: toneL = `g;     15'd367: toneL = `g;
                    // 15'd368: toneL = `g;     15'd369: toneL = `g;
                    // 15'd370: toneL = `g;     15'd371: toneL = `g;
                    // 15'd372: toneL = `g;     15'd373: toneL = `g;
                    // 15'd374: toneL = `g;     15'd375: toneL = `g;
                    // 15'd376: toneL = `sil;     15'd377: toneL = `sil;
                    // 15'd378: toneL = `g;     15'd379: toneL = `g;
                    // 15'd380: toneL = `g;     15'd381: toneL = `g;
                    // 15'd382: toneL = `g;     15'd383: toneL = `g;
                    // 15'd384: toneL = `g;     15'd385: toneL = `g;
                    // 15'd386: toneL = `g;     15'd387: toneL = `g;
                    // 15'd388: toneL = `g;     15'd389: toneL = `g;
                    // 15'd390: toneL = `g;     15'd391: toneL = `g;
                    // 15'd392: toneL = `g;     15'd393: toneL = `g;
                    // 15'd394: toneL = `g;     15'd395: toneL = `g;
                    // 15'd396: toneL = `g;     15'd397: toneL = `g;
                    // 15'd398: toneL = `g;     15'd399: toneL = `g;
                    // 15'd400: toneL = `g;     15'd401: toneL = `g;
                    // 15'd402: toneL = `g;     15'd403: toneL = `g;
                    // 15'd404: toneL = `g;     15'd405: toneL = `g;
                    // 15'd406: toneL = `g;     15'd407: toneL = `g;
                    // 15'd408: toneL = `g;     15'd409: toneL = `g;
                    // 15'd410: toneL = `g;     15'd411: toneL = `g;
                    // 15'd412: toneL = `g;     15'd413: toneL = `g;
                    // 15'd414: toneL = `g;     15'd415: toneL = `g;
                    // 15'd416: toneL = `e;     15'd417: toneL = `e;
                    // 15'd418: toneL = `e;     15'd419: toneL = `e;
                    // 15'd420: toneL = `e;     15'd421: toneL = `e;
                    // 15'd422: toneL = `e;     15'd423: toneL = `e;
                    // 15'd424: toneL = `e;     15'd425: toneL = `e;
                    // 15'd426: toneL = `e;     15'd427: toneL = `e;
                    // 15'd428: toneL = `e;     15'd429: toneL = `e;
                    // 15'd430: toneL = `e;     15'd431: toneL = `e;
                    // 15'd432: toneL = `e;     15'd433: toneL = `e;
                    // 15'd434: toneL = `e;     15'd435: toneL = `e;
                    // 15'd436: toneL = `e;     15'd437: toneL = `e;
                    // 15'd438: toneL = `e;     15'd439: toneL = `e;
                    // 15'd440: toneL = `e;     15'd441: toneL = `e;
                    // 15'd442: toneL = `e;     15'd443: toneL = `e;
                    // 15'd444: toneL = `e;     15'd445: toneL = `e;
                    // 15'd446: toneL = `e;     15'd447: toneL = `e;
                    // 15'd448: toneL = `g;     15'd449: toneL = `g;
                    // 15'd450: toneL = `g;     15'd451: toneL = `g;
                    // 15'd452: toneL = `g;     15'd453: toneL = `g;
                    // 15'd454: toneL = `g;     15'd455: toneL = `g;
                    // 15'd456: toneL = `g;     15'd457: toneL = `g;
                    // 15'd458: toneL = `g;     15'd459: toneL = `g;
                    // 15'd460: toneL = `g;     15'd461: toneL = `g;
                    // 15'd462: toneL = `g;     15'd463: toneL = `g;
                    // 15'd464: toneL = `g;     15'd465: toneL = `g;
                    // 15'd466: toneL = `g;     15'd467: toneL = `g;
                    // 15'd468: toneL = `g;     15'd469: toneL = `g;
                    // 15'd470: toneL = `g;     15'd471: toneL = `g;
                    // 15'd472: toneL = `g;     15'd473: toneL = `g;
                    // 15'd474: toneL = `g;     15'd475: toneL = `g;
                    // 15'd476: toneL = `g;     15'd477: toneL = `g;
                    // 15'd478: toneL = `g;     15'd479: toneL = `g;
                    // 15'd480: toneL = `e;     15'd481: toneL = `e;
                    // 15'd482: toneL = `e;     15'd483: toneL = `e;
                    // 15'd484: toneL = `e;     15'd485: toneL = `e;
                    // 15'd486: toneL = `e;     15'd487: toneL = `e;
                    // 15'd488: toneL = `e;     15'd489: toneL = `e;
                    // 15'd490: toneL = `e;     15'd491: toneL = `e;
                    // 15'd492: toneL = `e;     15'd493: toneL = `e;
                    // 15'd494: toneL = `e;     15'd495: toneL = `e;
                    // 15'd496: toneL = `e;     15'd497: toneL = `e;
                    // 15'd498: toneL = `e;     15'd499: toneL = `e;
                    // 15'd500: toneL = `e;     15'd501: toneL = `e;
                    // 15'd502: toneL = `e;     15'd503: toneL = `e;
                    // 15'd504: toneL = `e;     15'd505: toneL = `e;
                    // 15'd506: toneL = `e;     15'd507: toneL = `e;
                    // 15'd508: toneL = `e;     15'd509: toneL = `e;
                    // 15'd510: toneL = `e;     15'd511: toneL = `e;
        //         default : toneL = `sil;
        //     endcase
        end
         else begin
             toneL = `sil;
         end
    end

    //  always @(*) begin
    //     if(en == 1) begin
    //         case(ibeatNum)
    //             12'd0: TONE = `GG;  	12'd1: TONE = `GG; // HC (two-beat)
    //             12'd2: TONE = `GG;  	12'd3: TONE = `GG;
    //             12'd4: TONE = `GG;	    12'd5: TONE = `GG;
    //             12'd6: TONE = `GG;  	12'd7: TONE = `GG;
    //             12'd8: TONE = `AA;	    12'd9: TONE = `AA;
    //             12'd10: TONE = `AA;	12'd11: TONE = `AA;
    //             12'd12: TONE = `AA;	12'd13: TONE = `AA;
    //             12'd14: TONE = `AA;	12'd15: TONE = `AA;

    //             12'd16: TONE = `AA;	12'd17: TONE = `AA;
    //             12'd18: TONE = `GG;	12'd19: TONE = `GG;
    //             12'd20: TONE = `GG;	12'd21: TONE = `GG;
    //             12'd22: TONE = `GG;	12'd23: TONE = `GG;
    //             12'd24: TONE = `GG;	12'd25: TONE = `GG;
    //             12'd26: TONE = `GG;	12'd27: TONE = `GG;
    //             12'd28: TONE = `GG;	12'd29: TONE = `GG;
    //             12'd30: TONE = `GG;	12'd31: TONE = `GG;
    //             default : TONE = `BB;
    //         endcase
    //     end
    //     else begin
    //         TONE = `sil;
    //     end
    // end
endmodule